magic
tech sky130A
magscale 1 2
timestamp 1757527180
<< viali >>
rect 6481 -1695 6656 -1661
rect 13369 -2552 13409 -2512
rect 8297 -2928 8338 -2894
rect 9070 -2937 9119 -2888
rect 9965 -2928 10047 -2894
rect 11388 -3256 11436 -3222
rect 12883 -3574 12919 -3540
rect 13285 -3579 13334 -3545
rect 9156 -3720 9196 -3680
rect 10188 -3910 10230 -3876
rect 6524 -3965 6667 -3931
rect 11388 -4039 11449 -4005
rect 11388 -4260 11449 -4226
rect 8260 -4332 8294 -4298
rect 6524 -4372 6667 -4338
rect 11562 -4714 11711 -4680
rect 7769 -4849 7820 -4798
rect 11562 -5000 11711 -4966
rect 11399 -5454 11535 -5420
rect 10074 -5726 10126 -5692
rect 8276 -5824 8310 -5790
rect 8324 -7064 8452 -7030
<< metal1 >>
rect 5970 -1330 6170 -1329
rect 5970 -1529 13792 -1330
rect 5971 -1530 6170 -1529
rect 6469 -1661 6668 -1529
rect 6469 -1695 6481 -1661
rect 6656 -1695 6668 -1661
rect 6469 -1772 6668 -1695
rect 6774 -2116 8601 -2050
rect 8667 -2116 8673 -2050
rect 6540 -2222 6592 -2216
rect 6540 -2280 6592 -2274
rect 9063 -2314 9115 -2308
rect 8130 -2344 8837 -2316
rect 8130 -2372 8162 -2344
rect 8809 -2383 8837 -2344
rect 9063 -2372 9115 -2366
rect 7647 -2589 8140 -2561
rect 5992 -2860 6374 -2753
rect 5992 -5375 6099 -2860
rect 8291 -2894 8344 -2818
rect 8291 -2928 8297 -2894
rect 8338 -2928 8344 -2894
rect 8291 -3033 8344 -2928
rect 6907 -3182 6942 -3054
rect 8343 -3085 8344 -3033
rect 8291 -3108 8344 -3085
rect 9064 -2888 9125 -2820
rect 9064 -2937 9070 -2888
rect 9119 -2929 9125 -2888
rect 9516 -2929 9577 -1529
rect 9990 -2314 10042 -2308
rect 9726 -2362 9805 -2316
rect 9726 -2372 9772 -2362
rect 9990 -2372 10042 -2366
rect 9119 -2937 9577 -2929
rect 9064 -2990 9577 -2937
rect 9064 -3108 9125 -2990
rect 9726 -3164 9760 -2720
rect 9959 -2894 10053 -2820
rect 9959 -2928 9965 -2894
rect 10047 -2928 10053 -2894
rect 9959 -2938 10053 -2928
rect 9959 -2990 10677 -2938
rect 9959 -3033 10053 -2990
rect 9959 -3085 9977 -3033
rect 10029 -3085 10053 -3033
rect 9959 -3108 10053 -3085
rect 6893 -3188 6957 -3182
rect 6893 -3240 6899 -3188
rect 6951 -3240 6957 -3188
rect 6893 -3246 6957 -3240
rect 6907 -3353 6942 -3246
rect 6167 -3624 6173 -3535
rect 6262 -3624 6384 -3535
rect 10625 -3536 10677 -2990
rect 11396 -3204 11432 -1529
rect 12432 -2633 12520 -1529
rect 13202 -2305 13268 -2249
rect 13422 -2506 13474 -1529
rect 13624 -2305 13690 -2249
rect 13302 -2512 13592 -2506
rect 13040 -2571 13172 -2517
rect 13302 -2552 13369 -2512
rect 13409 -2552 13592 -2512
rect 13302 -2558 13592 -2552
rect 11376 -3222 11449 -3204
rect 11376 -3256 11388 -3222
rect 11436 -3256 11449 -3222
rect 11376 -3270 11449 -3256
rect 11690 -3262 11696 -3210
rect 11748 -3217 11754 -3210
rect 11748 -3254 12126 -3217
rect 11748 -3262 11754 -3254
rect 13040 -3284 13094 -2571
rect 13713 -2596 13882 -2542
rect 13936 -2596 13942 -2542
rect 13208 -2787 13262 -2786
rect 13202 -2792 13268 -2787
rect 13202 -2846 13208 -2792
rect 13262 -2803 13268 -2792
rect 13262 -2846 13333 -2803
rect 13624 -2806 13690 -2787
rect 13882 -2792 13936 -2596
rect 13202 -2859 13333 -2846
rect 13277 -3117 13333 -2859
rect 13623 -2862 13755 -2806
rect 13699 -3117 13755 -2862
rect 13936 -2846 13942 -2792
rect 13277 -3173 13343 -3117
rect 13699 -3173 13765 -3117
rect 13882 -3226 13936 -2846
rect 13797 -3280 13936 -3226
rect 11004 -3322 11056 -3316
rect 11376 -3321 11428 -3315
rect 11004 -3380 11056 -3374
rect 8132 -3584 8160 -3555
rect 8805 -3556 8830 -3541
rect 8805 -3584 8833 -3556
rect 8132 -3612 8833 -3584
rect 9292 -3612 9808 -3584
rect 10625 -3594 10677 -3588
rect 8132 -3829 8160 -3612
rect 9144 -3726 9150 -3674
rect 9202 -3726 9208 -3674
rect 7647 -3857 8160 -3829
rect 9558 -3798 9586 -3612
rect 10946 -3666 10952 -3607
rect 9558 -3826 10854 -3798
rect 6516 -3931 6673 -3915
rect 6516 -3965 6524 -3931
rect 6667 -3965 6673 -3931
rect 6516 -4338 6673 -3965
rect 9558 -4144 9586 -3826
rect 10170 -3876 10248 -3863
rect 10170 -3910 10188 -3876
rect 10230 -3910 10248 -3876
rect 10170 -3923 10248 -3910
rect 10170 -3975 10189 -3923
rect 10241 -3975 10248 -3923
rect 10170 -3984 10248 -3975
rect 9558 -4172 9930 -4144
rect 6516 -4372 6524 -4338
rect 6667 -4342 6673 -4338
rect 8254 -4298 8300 -4286
rect 8254 -4332 8260 -4298
rect 8294 -4332 8300 -4298
rect 6667 -4370 7238 -4342
rect 8254 -4344 8300 -4332
rect 6667 -4372 6673 -4370
rect 6516 -4386 6673 -4372
rect 6562 -4446 6627 -4386
rect 7210 -4475 7238 -4370
rect 8263 -4405 8291 -4344
rect 10826 -4390 10854 -3826
rect 11011 -3883 11048 -3380
rect 11246 -3430 11302 -3364
rect 11376 -3379 11428 -3373
rect 11514 -3367 11570 -3364
rect 11514 -3421 11939 -3367
rect 11993 -3421 11999 -3367
rect 11514 -3430 11570 -3421
rect 11388 -3624 11447 -3464
rect 12688 -3467 12723 -3334
rect 13094 -3338 13245 -3284
rect 13377 -3338 13667 -3286
rect 13040 -3344 13094 -3338
rect 12688 -3502 13200 -3467
rect 13277 -3493 13343 -3437
rect 12688 -3563 12723 -3502
rect 12875 -3538 12927 -3532
rect 11995 -3598 12723 -3563
rect 12871 -3575 12875 -3540
rect 12927 -3575 12931 -3540
rect 12875 -3596 12927 -3590
rect 11995 -3624 12030 -3598
rect 11388 -3659 12030 -3624
rect 12688 -3648 12723 -3598
rect 11388 -3797 11447 -3659
rect 11004 -3889 11056 -3883
rect 11288 -3897 11344 -3831
rect 11492 -3836 11548 -3831
rect 11384 -3888 11436 -3882
rect 11004 -3947 11056 -3941
rect 11492 -3890 12306 -3836
rect 12360 -3890 12366 -3836
rect 11492 -3897 11548 -3890
rect 11384 -3946 11436 -3940
rect 11376 -4005 11460 -3994
rect 11376 -4039 11388 -4005
rect 11449 -4039 11461 -4005
rect 11376 -4226 11461 -4039
rect 11956 -4045 11962 -3993
rect 12014 -4000 12020 -3993
rect 12014 -4037 12612 -4000
rect 12014 -4045 12020 -4037
rect 11376 -4260 11388 -4226
rect 11449 -4260 11461 -4226
rect 11376 -4273 11461 -4260
rect 12758 -4323 12810 -4317
rect 12758 -4381 12810 -4375
rect 8261 -4433 8933 -4405
rect 10826 -4418 10862 -4390
rect 8543 -4667 8848 -4631
rect 10099 -4791 10165 -4488
rect 11613 -4671 11677 -4618
rect 11613 -4674 11619 -4671
rect 11550 -4680 11619 -4674
rect 11671 -4674 11677 -4671
rect 11671 -4680 11723 -4674
rect 11550 -4714 11562 -4680
rect 11711 -4714 11723 -4680
rect 11550 -4720 11619 -4714
rect 11613 -4723 11619 -4720
rect 11671 -4720 11723 -4714
rect 11671 -4723 11677 -4720
rect 12302 -4791 12330 -4540
rect 13165 -4791 13200 -3502
rect 13284 -3533 13336 -3532
rect 13279 -3535 13340 -3533
rect 13496 -3535 13548 -3338
rect 13279 -3538 13548 -3535
rect 13279 -3590 13284 -3538
rect 13336 -3587 13548 -3538
rect 13699 -3493 13765 -3437
rect 13336 -3590 13340 -3587
rect 13279 -3591 13340 -3590
rect 13284 -3596 13336 -3591
rect 13699 -3700 13756 -3493
rect 13805 -3700 14005 -3629
rect 13699 -3757 14005 -3700
rect 13805 -3829 14005 -3757
rect 13805 -4791 14005 -4666
rect 7757 -4855 7763 -4792
rect 7826 -4855 7832 -4792
rect 8285 -4863 8337 -4857
rect 8518 -4863 8564 -4847
rect 6888 -4903 6934 -4870
rect 6642 -5248 6670 -4933
rect 6847 -4950 6934 -4903
rect 6887 -5097 6934 -4950
rect 7171 -4918 7223 -4912
rect 7668 -4916 7714 -4875
rect 7223 -4958 7286 -4930
rect 7640 -4962 7714 -4916
rect 8477 -4909 8564 -4863
rect 10099 -4857 14005 -4791
rect 8285 -4921 8337 -4915
rect 7171 -4976 7223 -4970
rect 6887 -5110 8027 -5097
rect 6888 -5144 8027 -5110
rect 7996 -5312 8027 -5144
rect 8930 -5211 8958 -4884
rect 10099 -5114 10165 -4857
rect 11613 -4959 11619 -4956
rect 11550 -4966 11619 -4959
rect 11671 -4959 11677 -4956
rect 11671 -4966 11723 -4959
rect 11550 -5000 11562 -4966
rect 11711 -5000 11723 -4966
rect 11550 -5006 11619 -5000
rect 11613 -5008 11619 -5006
rect 11671 -5006 11723 -5000
rect 11671 -5008 11677 -5006
rect 11613 -5062 11677 -5008
rect 12302 -5147 12330 -4857
rect 13805 -4866 14005 -4857
rect 8474 -5239 9936 -5211
rect 10279 -5249 10830 -5198
rect 8848 -5292 8900 -5286
rect 8848 -5350 8900 -5344
rect 5945 -5428 6145 -5375
rect 5945 -5521 6381 -5428
rect 7763 -5432 7826 -5426
rect 5945 -5575 6145 -5521
rect 6600 -6048 6631 -5718
rect 6821 -5742 7083 -5714
rect 5945 -6231 6145 -6176
rect 5945 -6320 6173 -6231
rect 6262 -6320 6362 -6231
rect 7055 -6244 7083 -5742
rect 7763 -5990 7826 -5495
rect 8275 -5784 8311 -5713
rect 8270 -5790 8316 -5784
rect 8270 -5824 8276 -5790
rect 8310 -5824 8316 -5790
rect 8270 -5830 8316 -5824
rect 8602 -5821 8654 -5815
rect 8275 -6244 8311 -5830
rect 8602 -5879 8654 -5873
rect 8614 -6007 8642 -5879
rect 8860 -6068 8888 -5350
rect 11387 -5420 11547 -5414
rect 11387 -5454 11399 -5420
rect 11535 -5454 11547 -5420
rect 11387 -5462 11547 -5454
rect 10074 -5685 10126 -5616
rect 10068 -5692 10132 -5685
rect 10068 -5726 10074 -5692
rect 10126 -5726 10132 -5692
rect 10068 -5732 10132 -5726
rect 10074 -5929 10126 -5732
rect 11454 -5929 11485 -5462
rect 10074 -5960 11485 -5929
rect 7055 -6272 7207 -6244
rect 8078 -6280 8407 -6244
rect 5945 -6376 6145 -6320
rect 6719 -6486 6771 -6480
rect 6719 -6544 6771 -6538
rect 8142 -6654 8194 -6648
rect 7955 -6691 8142 -6663
rect 5945 -6856 6145 -6770
rect 7955 -6824 7983 -6691
rect 8194 -6691 8329 -6663
rect 8142 -6712 8194 -6706
rect 8301 -6827 8329 -6691
rect 5945 -6922 6406 -6856
rect 8070 -6922 8224 -6855
rect 9888 -6922 9944 -6856
rect 5945 -6970 6145 -6922
rect 7533 -7143 7561 -6939
rect 8312 -7030 8464 -7024
rect 8312 -7064 8324 -7030
rect 8452 -7064 8464 -7030
rect 8312 -7086 8464 -7064
rect 8381 -7143 8409 -7086
rect 8775 -7143 8803 -6948
rect 7533 -7171 8803 -7143
rect 8137 -7289 8165 -7171
rect 10074 -7289 10126 -5960
rect 11799 -7224 11805 -7159
rect 11870 -7224 11876 -7159
rect 11805 -7289 11870 -7224
rect 5945 -7489 12033 -7289
<< via1 >>
rect 8601 -2116 8667 -2050
rect 6540 -2274 6592 -2222
rect 9063 -2366 9115 -2314
rect 8291 -3085 8343 -3033
rect 9990 -2366 10042 -2314
rect 9977 -3085 10029 -3033
rect 6899 -3240 6951 -3188
rect 6173 -3624 6262 -3535
rect 11696 -3262 11748 -3210
rect 13882 -2596 13936 -2542
rect 13208 -2846 13262 -2792
rect 13882 -2846 13936 -2792
rect 11004 -3374 11056 -3322
rect 10625 -3588 10677 -3536
rect 9150 -3680 9202 -3674
rect 9150 -3720 9156 -3680
rect 9156 -3720 9196 -3680
rect 9196 -3720 9202 -3680
rect 9150 -3726 9202 -3720
rect 10952 -3666 11011 -3607
rect 10189 -3975 10241 -3923
rect 11376 -3373 11428 -3321
rect 11939 -3421 11993 -3367
rect 13040 -3338 13094 -3284
rect 12875 -3540 12927 -3538
rect 12875 -3574 12883 -3540
rect 12883 -3574 12919 -3540
rect 12919 -3574 12927 -3540
rect 12875 -3590 12927 -3574
rect 11004 -3941 11056 -3889
rect 11384 -3940 11436 -3888
rect 12306 -3890 12360 -3836
rect 11962 -4045 12014 -3993
rect 12758 -4375 12810 -4323
rect 11619 -4680 11671 -4671
rect 11619 -4714 11671 -4680
rect 11619 -4723 11671 -4714
rect 13284 -3545 13336 -3538
rect 13284 -3579 13285 -3545
rect 13285 -3579 13334 -3545
rect 13334 -3579 13336 -3545
rect 13284 -3590 13336 -3579
rect 7763 -4798 7826 -4792
rect 7763 -4849 7769 -4798
rect 7769 -4849 7820 -4798
rect 7820 -4849 7826 -4798
rect 7763 -4855 7826 -4849
rect 7171 -4970 7223 -4918
rect 8285 -4915 8337 -4863
rect 11619 -4966 11671 -4956
rect 11619 -5000 11671 -4966
rect 11619 -5008 11671 -5000
rect 8848 -5344 8900 -5292
rect 7763 -5495 7826 -5432
rect 6173 -6320 6262 -6231
rect 8602 -5873 8654 -5821
rect 6719 -6538 6771 -6486
rect 8142 -6706 8194 -6654
rect 11805 -7224 11870 -7159
<< metal2 >>
rect 8601 -2050 8667 -2044
rect 6534 -2274 6540 -2222
rect 6592 -2231 6598 -2222
rect 6592 -2266 7825 -2231
rect 6592 -2274 6598 -2266
rect 6893 -3188 6957 -3182
rect 6893 -3240 6899 -3188
rect 6951 -3196 6957 -3188
rect 7790 -3196 7825 -2266
rect 8601 -3033 8667 -2116
rect 11939 -2210 13936 -2156
rect 9057 -2366 9063 -2314
rect 9115 -2326 9121 -2314
rect 9984 -2326 9990 -2314
rect 9115 -2354 9990 -2326
rect 9115 -2366 9121 -2354
rect 9984 -2366 9990 -2354
rect 10042 -2366 10048 -2314
rect 8285 -3085 8291 -3033
rect 8343 -3085 9977 -3033
rect 10029 -3085 10035 -3033
rect 6951 -3231 7825 -3196
rect 11696 -3210 11748 -3204
rect 6951 -3240 6957 -3231
rect 6893 -3246 6957 -3240
rect 11696 -3268 11748 -3262
rect 10998 -3374 11004 -3322
rect 11056 -3329 11062 -3322
rect 11370 -3329 11376 -3321
rect 11056 -3366 11376 -3329
rect 11056 -3374 11062 -3366
rect 11370 -3373 11376 -3366
rect 11428 -3329 11434 -3321
rect 11703 -3329 11740 -3268
rect 11428 -3366 11740 -3329
rect 11428 -3373 11434 -3366
rect 11939 -3367 11993 -2210
rect 13882 -2542 13936 -2210
rect 13882 -2602 13936 -2596
rect 13202 -2846 13208 -2792
rect 13262 -2846 13882 -2792
rect 13936 -2846 13942 -2792
rect 13034 -3338 13040 -3284
rect 13094 -3338 13100 -3284
rect 13040 -3371 13094 -3338
rect 11939 -3427 11993 -3421
rect 12306 -3425 13094 -3371
rect 10952 -3449 11012 -3440
rect 10952 -3518 11012 -3509
rect 6173 -3535 6262 -3529
rect 10619 -3588 10625 -3536
rect 10677 -3588 10683 -3536
rect 6173 -6231 6262 -3624
rect 9150 -3674 9202 -3668
rect 9150 -3732 9202 -3726
rect 9160 -3936 9191 -3732
rect 10189 -3923 10241 -3917
rect 9160 -3967 10189 -3936
rect 10189 -3981 10241 -3975
rect 10625 -4672 10677 -3588
rect 10952 -3607 11011 -3518
rect 10952 -3672 11011 -3666
rect 12306 -3836 12360 -3425
rect 12869 -3590 12875 -3538
rect 12927 -3550 12933 -3538
rect 13278 -3550 13284 -3538
rect 12927 -3578 13284 -3550
rect 12927 -3590 12933 -3578
rect 13278 -3590 13284 -3578
rect 13336 -3590 13342 -3538
rect 10998 -3941 11004 -3889
rect 11056 -3896 11062 -3889
rect 11378 -3896 11384 -3888
rect 11056 -3933 11384 -3896
rect 11056 -3941 11062 -3933
rect 11378 -3940 11384 -3933
rect 11436 -3896 11442 -3888
rect 12306 -3896 12360 -3890
rect 11436 -3933 12006 -3896
rect 11436 -3940 11442 -3933
rect 11969 -3987 12006 -3933
rect 11962 -3993 12014 -3987
rect 11962 -4051 12014 -4045
rect 12752 -4375 12758 -4323
rect 12810 -4375 12816 -4323
rect 11619 -4671 11671 -4665
rect 10625 -4723 11619 -4672
rect 10625 -4724 11671 -4723
rect 11619 -4729 11671 -4724
rect 7763 -4792 7826 -4786
rect 7165 -4930 7171 -4918
rect 6173 -6326 6262 -6320
rect 7012 -4958 7171 -4930
rect 7012 -5833 7040 -4958
rect 7165 -4970 7171 -4958
rect 7223 -4970 7229 -4918
rect 7763 -5432 7826 -4855
rect 8279 -4915 8285 -4863
rect 8337 -4875 8343 -4863
rect 8337 -4903 8888 -4875
rect 8337 -4915 8343 -4903
rect 8860 -5292 8888 -4903
rect 11631 -4950 11659 -4729
rect 11619 -4956 11671 -4950
rect 11619 -5014 11671 -5008
rect 8842 -5344 8848 -5292
rect 8900 -5344 8906 -5292
rect 7757 -5495 7763 -5432
rect 7826 -5495 7832 -5432
rect 8596 -5833 8602 -5821
rect 7012 -5861 8602 -5833
rect 6713 -6538 6719 -6486
rect 6771 -6498 6777 -6486
rect 7012 -6498 7040 -5861
rect 8596 -5873 8602 -5861
rect 8654 -5873 8660 -5821
rect 6771 -6526 7040 -6498
rect 6771 -6538 6777 -6526
rect 8136 -6706 8142 -6654
rect 8194 -6666 8200 -6654
rect 12770 -6666 12798 -4375
rect 8194 -6694 12798 -6666
rect 8194 -6706 8200 -6694
rect 11805 -6991 11870 -6986
rect 11800 -7047 11809 -6991
rect 11865 -7047 11874 -6991
rect 11805 -7159 11870 -7047
rect 11805 -7230 11870 -7224
<< via2 >>
rect 10952 -3509 11012 -3449
rect 11809 -7047 11865 -6991
<< metal3 >>
rect 10950 -3286 11014 -3280
rect 10950 -3356 11014 -3350
rect 10952 -3444 11012 -3356
rect 10947 -3449 11017 -3444
rect 10947 -3509 10952 -3449
rect 11012 -3509 11017 -3449
rect 10947 -3514 11017 -3509
rect 11804 -6823 11869 -6822
rect 11798 -6887 11804 -6823
rect 11868 -6887 11874 -6823
rect 11804 -6986 11869 -6887
rect 11804 -6991 11870 -6986
rect 11804 -7047 11809 -6991
rect 11865 -7047 11870 -6991
rect 11804 -7052 11870 -7047
<< via3 >>
rect 10950 -3350 11014 -3286
rect 11804 -6887 11868 -6823
<< metal4 >>
rect 10952 -3285 11012 -3055
rect 10949 -3286 11015 -3285
rect 10949 -3350 10950 -3286
rect 11014 -3350 11015 -3286
rect 10949 -3351 11015 -3350
rect 11803 -6822 11868 -3091
rect 11803 -6823 11869 -6822
rect 11803 -6887 11804 -6823
rect 11868 -6887 11869 -6823
rect 11803 -6888 11869 -6887
use sky130_fd_pr__cap_mim_m3_1_BZXCPH  XC4
timestamp 1757456334
transform 1 0 11304 0 1 -2598
box -586 -540 586 540
use sky130_fd_pr__nfet_01v8_XVWV9Z  XM1
timestamp 1757456334
transform 0 1 6639 -1 0 -6282
box -396 -410 396 410
use sky130_fd_pr__nfet_01v8_XVWV9Z  XM2
timestamp 1757456334
transform 0 1 6638 -1 0 -5490
box -396 -410 396 410
use sky130_fd_pr__nfet_01v8_FMZK9W  XM3
timestamp 1757456334
transform 1 0 7645 0 1 -6268
box -596 -410 596 410
use sky130_fd_pr__pfet_01v8_lvt_GW5SVV  XM4
timestamp 1757456334
transform -1 0 7462 0 -1 -4675
box -396 -419 396 419
use sky130_fd_pr__pfet_01v8_lvt_GW5SVV  XM5
timestamp 1757456334
transform 0 1 6647 -1 0 -4697
box -396 -419 396 419
use sky130_fd_pr__pfet_01v8_GJP7VV  XM6
timestamp 1757456334
transform 0 1 7047 -1 0 -3605
box -396 -819 396 819
use sky130_fd_pr__pfet_01v8_GJP7VV  XM7
timestamp 1757456334
transform 0 1 7047 -1 0 -2813
box -396 -819 396 819
use sky130_fd_pr__nfet_01v8_lvt_L3FTKF  XM8
timestamp 1757456334
transform 0 1 8310 -1 0 -3360
box -396 -310 396 310
use sky130_fd_pr__nfet_01v8_lvt_L3FTKF  XM9
timestamp 1757456334
transform 0 1 8308 -1 0 -2568
box -396 -310 396 310
use sky130_fd_pr__pfet_01v8_8JYSVV  XM10
timestamp 1757456334
transform 0 1 6567 -1 0 -2021
box -396 -339 396 339
use sky130_fd_pr__nfet_01v8_lvt_XVWV9Z  XM11
timestamp 1757456334
transform 1 0 8636 0 1 -6266
box -396 -410 396 410
use sky130_fd_pr__nfet_01v8_lvt_XVWV9Z  XM12
timestamp 1757456334
transform 0 1 8274 -1 0 -5463
box -396 -410 396 410
use sky130_fd_pr__pfet_01v8_lvt_GW5SVV  XM13
timestamp 1757456334
transform 0 1 8277 -1 0 -4658
box -396 -419 396 419
use sky130_fd_pr__pfet_01v8_lvt_GW5SVV  XM14
timestamp 1757456334
transform 0 1 9115 -1 0 -4658
box -396 -419 396 419
use sky130_fd_pr__nfet_01v8_lvt_XVWV9Z  XM15
timestamp 1757456334
transform 0 1 10004 -1 0 -3360
box -396 -410 396 410
use sky130_fd_pr__nfet_01v8_lvt_XVWV9Z  XM16
timestamp 1757456334
transform 0 1 10004 -1 0 -2568
box -396 -410 396 410
use sky130_fd_pr__pfet_01v8_lvt_GW5SVV  XM17
timestamp 1757456334
transform 0 1 9096 -1 0 -2568
box -396 -419 396 419
use sky130_fd_pr__pfet_01v8_lvt_GW5SVV  XM18
timestamp 1757456334
transform 0 1 9096 -1 0 -3360
box -396 -419 396 419
use sky130_fd_pr__nfet_01v8_L3FTKF  XM19
timestamp 1757456334
transform 0 1 10101 -1 0 -5366
box -396 -310 396 310
use sky130_fd_pr__pfet_01v8_GJB8VV  XM20
timestamp 1757456334
transform 0 1 10207 -1 0 -4236
box -396 -419 396 419
use sky130_fd_pr__nfet_01v8_FMD5LY  XM21
timestamp 1757456334
transform 1 0 11578 0 1 -5210
box -896 -280 896 280
use sky130_fd_pr__nfet_01v8_FMD5LY  XM22
timestamp 1757456334
transform 1 0 11578 0 1 -4470
box -896 -280 896 280
use sky130_fd_pr__nfet_01v8_lvt_V433WY  XM23
timestamp 1757456334
transform 0 1 12784 -1 0 -4000
box -496 -310 496 310
use sky130_fd_pr__pfet_01v8_lvt_CEYSV5  XM24
timestamp 1757456334
transform 0 1 12505 -1 0 -2985
box -496 -519 496 519
use sky130_fd_pr__pfet_01v8_XGAKDL  XM25
timestamp 1757456334
transform -1 0 13657 0 -1 -2546
box -211 -419 211 419
use sky130_fd_pr__nfet_01v8_648S5X  XM26
timestamp 1757456334
transform 1 0 13732 0 1 -3303
box -211 -310 211 310
use sky130_fd_pr__nfet_01v8_648S5X  XM27
timestamp 1757456334
transform 1 0 13310 0 1 -3305
box -211 -310 211 310
use sky130_fd_pr__pfet_01v8_XGAKDL  XM28
timestamp 1757456334
transform 1 0 13235 0 1 -2546
box -211 -419 211 419
use sky130_fd_pr__nfet_01v8_PWNS5P  XM29
timestamp 1757456334
transform 0 1 8147 -1 0 -6889
box -211 -1919 211 1919
use sky130_fd_pr__pfet_01v8_X6BGBL  XM30
timestamp 1757456334
transform 0 1 11413 -1 0 -3397
box -211 -289 211 289
use sky130_fd_pr__nfet_01v8_L7T3GD  XM31
timestamp 1757456334
transform 0 1 11418 -1 0 -3864
box -211 -252 211 252
<< labels >>
flabel metal1 8930 -5239 8958 -4884 0 FreeSans 160 0 0 0 out2
flabel space 9280 -3612 9816 -3584 0 FreeSans 320 0 0 0 out1
flabel space 11011 -3666 12150 -3607 0 FreeSans 320 0 0 0 ZERO0
flabel metal1 5945 -6970 6145 -6770 0 FreeSans 256 0 0 0 EN_N
port 0 nsew
flabel metal1 5945 -7489 6145 -7289 0 FreeSans 256 0 0 0 VSS
port 6 nsew
flabel metal1 5945 -6376 6145 -6176 0 FreeSans 256 0 0 0 PLUS
port 1 nsew
flabel metal1 13805 -4866 14005 -4666 0 FreeSans 256 0 0 0 comp_out
port 4 nsew
flabel metal1 13805 -3829 14005 -3629 0 FreeSans 256 0 0 0 CAL
port 3 nsew
flabel metal1 13882 -3280 13936 -2846 0 FreeSans 320 0 0 0 CALB
flabel metal1 13040 -3338 13094 -2517 0 FreeSans 320 0 0 0 CALBB
flabel metal1 7955 -6691 8329 -6663 0 FreeSans 320 0 0 0 VSSI
flabel metal1 11011 -3889 11025 -3885 0 FreeSans 320 0 0 0 ZERO0
flabel metal1 5945 -5575 6145 -5375 0 FreeSans 256 0 0 0 MINUS
port 2 nsew
flabel metal1 5970 -1529 6170 -1329 0 FreeSans 256 0 0 0 VCC
port 5 nsew
<< end >>
