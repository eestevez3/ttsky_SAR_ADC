** sch_path: /home/ttuser/ttsky_SAR_ADC/xschem/r2r_dac.sch
.subckt r2r_dac dac_out VSS b1 b3 b4 b5 b7 b6 b2 b0 VSUBS
*.PININFO b0:I dac_out:O b1:I b2:I b3:I b4:I b5:I b6:I b7:I VSS:I VSUBS:I
XR1 b0 dac_out VSUBS sky130_fd_pr__res_high_po_0p35 L=20 mult=1 m=1
XR2 dac_out net1 VSUBS sky130_fd_pr__res_high_po_0p35 L=10 mult=1 m=1
XR3 b1 net1 VSUBS sky130_fd_pr__res_high_po_0p35 L=20 mult=1 m=1
XR4 net1 net2 VSUBS sky130_fd_pr__res_high_po_0p35 L=10 mult=1 m=1
XR5 b2 net2 VSUBS sky130_fd_pr__res_high_po_0p35 L=20 mult=1 m=1
XR6 net2 net3 VSUBS sky130_fd_pr__res_high_po_0p35 L=10 mult=1 m=1
XR7 b3 net3 VSUBS sky130_fd_pr__res_high_po_0p35 L=20 mult=1 m=1
XR8 net3 net4 VSUBS sky130_fd_pr__res_high_po_0p35 L=10 mult=1 m=1
XR9 b4 net4 VSUBS sky130_fd_pr__res_high_po_0p35 L=20 mult=1 m=1
XR10 net4 net5 VSUBS sky130_fd_pr__res_high_po_0p35 L=10 mult=1 m=1
XR11 b5 net5 VSUBS sky130_fd_pr__res_high_po_0p35 L=20 mult=1 m=1
XR12 net5 net6 VSUBS sky130_fd_pr__res_high_po_0p35 L=10 mult=1 m=1
XR13 b6 net6 VSUBS sky130_fd_pr__res_high_po_0p35 L=20 mult=1 m=1
XR14 net6 net7 VSUBS sky130_fd_pr__res_high_po_0p35 L=10 mult=1 m=1
XR15 b7 net7 VSUBS sky130_fd_pr__res_high_po_0p35 L=20 mult=1 m=1
XR16 net7 VSS VSUBS sky130_fd_pr__res_high_po_0p35 L=20 mult=1 m=1
.ends
.end
