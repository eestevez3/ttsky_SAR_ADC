magic
tech sky130A
magscale 1 2
timestamp 1757456334
<< metal3 >>
rect -586 512 586 540
rect -586 -512 502 512
rect 566 -512 586 512
rect -586 -540 586 -512
<< via3 >>
rect 502 -512 566 512
<< mimcap >>
rect -546 460 254 500
rect -546 -460 -506 460
rect 214 -460 254 460
rect -546 -500 254 -460
<< mimcapcontact >>
rect -506 -460 214 460
<< metal4 >>
rect 486 512 582 528
rect -507 460 215 461
rect -507 -460 -506 460
rect 214 -460 215 460
rect -507 -461 215 -460
rect 486 -512 502 512
rect 566 -512 582 512
rect 486 -528 582 -512
<< properties >>
string FIXED_BBOX -586 -540 294 540
string gencell sky130_fd_pr__cap_mim_m3_1
string library sky130
string parameters w 4.0 l 5.0 val 43.42 carea 2.00 cperi 0.19 nx 1 ny 1 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1 ccov 100
<< end >>
