magic
tech sky130A
magscale 1 2
timestamp 1755657154
<< pwell >>
rect 727 -4230 911 -4225
rect 2822 -4229 2868 -4160
rect 1721 -4285 1905 -4230
rect 2706 -4284 2892 -4229
<< viali >>
rect 742 -3002 1004 -2968
rect 1736 -3002 1998 -2968
rect 2617 -3003 2879 -2969
rect 1640 -3339 1674 -3163
rect 2060 -3339 2094 -3163
rect 2521 -3340 2555 -3164
rect 2941 -3340 2975 -3164
rect 742 -4272 900 -4238
rect 1733 -4273 1891 -4239
rect 2722 -4272 2880 -4238
<< metal1 >>
rect 427 -2830 2891 -2630
rect 730 -2900 2891 -2830
rect 730 -2955 1015 -2900
rect 730 -2968 1016 -2955
rect 730 -3002 742 -2968
rect 1004 -3002 1016 -2968
rect 730 -3015 1016 -3002
rect 1725 -2968 2006 -2900
rect 1725 -3002 1736 -2968
rect 1998 -3002 2006 -2968
rect 1725 -3014 2006 -3002
rect 2605 -2969 2891 -2900
rect 2605 -3003 2617 -2969
rect 2879 -3003 2891 -2969
rect 2605 -3014 2891 -3003
rect 428 -3113 628 -3043
rect 885 -3110 1225 -3065
rect 428 -3172 627 -3113
rect 686 -3172 692 -3113
rect 428 -3243 628 -3172
rect 840 -3206 906 -3201
rect 740 -3258 746 -3206
rect 798 -3258 804 -3206
rect 840 -3258 848 -3206
rect 900 -3258 906 -3206
rect 840 -3265 906 -3258
rect 946 -3259 952 -3207
rect 1004 -3259 1010 -3207
rect 1180 -3225 1225 -3110
rect 1451 -3109 2207 -3064
rect 1451 -3112 1523 -3109
rect 1451 -3172 1457 -3112
rect 1517 -3172 1523 -3112
rect 1451 -3179 1523 -3172
rect 1628 -3163 1794 -3151
rect 1180 -3287 1301 -3225
rect 1363 -3287 1369 -3225
rect 1180 -3395 1225 -3287
rect 1628 -3339 1640 -3163
rect 1674 -3339 1794 -3163
rect 1940 -3163 2106 -3150
rect 1832 -3217 1896 -3211
rect 1832 -3269 1838 -3217
rect 1890 -3269 1896 -3217
rect 1832 -3275 1896 -3269
rect 1628 -3352 1794 -3339
rect 1940 -3339 2060 -3163
rect 2094 -3339 2106 -3163
rect 1940 -3351 2106 -3339
rect 2162 -3394 2207 -3109
rect 2377 -3109 2840 -3064
rect 785 -3440 1227 -3395
rect 1779 -3439 2207 -3394
rect 2162 -3496 2207 -3439
rect 2265 -3442 2271 -3390
rect 2323 -3394 2329 -3390
rect 2377 -3394 2422 -3109
rect 2509 -3164 2676 -3150
rect 2509 -3340 2521 -3164
rect 2555 -3340 2676 -3164
rect 2821 -3164 2988 -3150
rect 2717 -3228 2781 -3222
rect 2717 -3280 2723 -3228
rect 2775 -3280 2781 -3228
rect 2717 -3286 2781 -3280
rect 2509 -3352 2676 -3340
rect 2821 -3340 2941 -3164
rect 2975 -3340 2988 -3164
rect 2821 -3352 2988 -3340
rect 2323 -3439 2740 -3394
rect 2323 -3442 2329 -3439
rect 3231 -3468 3283 -3462
rect 2159 -3502 2211 -3496
rect 423 -3615 623 -3540
rect 3231 -3526 3283 -3520
rect 2159 -3560 2211 -3554
rect 952 -3614 1004 -3608
rect 2992 -3614 3192 -3537
rect 3231 -3614 3282 -3526
rect 423 -3667 746 -3615
rect 798 -3667 804 -3615
rect 1004 -3665 3282 -3614
rect 423 -3740 623 -3667
rect 952 -3672 1004 -3666
rect 2154 -3721 2160 -3718
rect 1793 -3766 2160 -3721
rect 1154 -3861 1229 -3856
rect 768 -3924 1160 -3861
rect 1223 -3924 1229 -3861
rect 1793 -3887 1838 -3766
rect 2154 -3770 2160 -3766
rect 2212 -3770 2218 -3718
rect 2992 -3737 3192 -3665
rect 783 -3928 862 -3924
rect 1154 -3932 1229 -3924
rect 1773 -3932 1853 -3887
rect 2114 -3932 2840 -3887
rect 740 -4079 746 -4027
rect 798 -4079 804 -4027
rect 842 -4085 848 -4033
rect 900 -4085 906 -4033
rect 1828 -4088 1834 -4026
rect 1896 -4046 1902 -4026
rect 2114 -4046 2159 -3932
rect 1896 -4088 2159 -4046
rect 2711 -4059 2717 -3996
rect 2780 -4059 2786 -3996
rect 1856 -4091 2159 -4088
rect 727 -4238 911 -4225
rect 1745 -4230 1791 -4120
rect 2822 -4229 2868 -4160
rect 727 -4272 742 -4238
rect 900 -4272 911 -4238
rect 727 -4391 911 -4272
rect 1721 -4239 1905 -4230
rect 1721 -4273 1733 -4239
rect 1891 -4273 1905 -4239
rect 1721 -4391 1905 -4273
rect 2706 -4238 2892 -4229
rect 2706 -4272 2722 -4238
rect 2880 -4272 2892 -4238
rect 2706 -4284 2892 -4272
rect 2706 -4391 2890 -4284
rect 727 -4405 2890 -4391
rect 424 -4494 2890 -4405
rect 424 -4598 3375 -4494
rect 3479 -4598 3485 -4494
rect 424 -4605 2890 -4598
<< via1 >>
rect 627 -3172 686 -3113
rect 746 -3258 798 -3206
rect 848 -3258 900 -3206
rect 952 -3259 1004 -3207
rect 1457 -3172 1517 -3112
rect 1301 -3287 1363 -3225
rect 1838 -3269 1890 -3217
rect 2271 -3442 2323 -3390
rect 2723 -3280 2775 -3228
rect 2159 -3554 2211 -3502
rect 3231 -3520 3283 -3468
rect 746 -3667 798 -3615
rect 952 -3666 1004 -3614
rect 1160 -3924 1223 -3861
rect 2160 -3770 2212 -3718
rect 746 -4079 798 -4027
rect 848 -4085 900 -4033
rect 1834 -4088 1896 -4026
rect 2717 -4059 2780 -3996
rect 3375 -4598 3479 -4494
<< metal2 >>
rect 619 -3112 696 -3102
rect 1459 -3106 1515 -3105
rect 619 -3172 627 -3112
rect 687 -3172 696 -3112
rect 1451 -3112 1524 -3106
rect 619 -3181 696 -3172
rect 758 -3150 992 -3122
rect 758 -3200 786 -3150
rect 746 -3206 798 -3200
rect 964 -3201 992 -3150
rect 1451 -3172 1457 -3112
rect 1517 -3172 1524 -3112
rect 1451 -3180 1524 -3172
rect 746 -3615 798 -3258
rect 840 -3206 906 -3201
rect 840 -3258 848 -3206
rect 900 -3258 906 -3206
rect 840 -3265 906 -3258
rect 952 -3207 1004 -3201
rect 1832 -3217 1896 -3211
rect 952 -3265 1004 -3259
rect 1301 -3225 1363 -3219
rect 746 -4027 798 -3667
rect 746 -4085 798 -4079
rect 848 -3615 899 -3265
rect 1832 -3269 1838 -3217
rect 1890 -3269 1896 -3217
rect 1832 -3275 1896 -3269
rect 946 -3615 952 -3614
rect 848 -3666 952 -3615
rect 1004 -3666 1010 -3614
rect 1301 -3651 1363 -3287
rect 1834 -3393 1896 -3275
rect 2717 -3228 2781 -3222
rect 2717 -3280 2723 -3228
rect 2775 -3280 2781 -3228
rect 2717 -3286 2781 -3280
rect 2271 -3390 2323 -3384
rect 1834 -3438 2271 -3393
rect 1834 -3651 1896 -3438
rect 2271 -3448 2323 -3442
rect 2153 -3554 2159 -3502
rect 2211 -3554 2217 -3502
rect 848 -4027 899 -3666
rect 1301 -3713 1896 -3651
rect 2163 -3712 2208 -3554
rect 2717 -3680 2780 -3286
rect 3228 -3310 3288 -3301
rect 3228 -3379 3288 -3370
rect 3232 -3468 3283 -3379
rect 3225 -3520 3231 -3468
rect 3283 -3520 3289 -3468
rect 1154 -3861 1229 -3856
rect 1154 -3924 1160 -3861
rect 1223 -3924 1229 -3861
rect 1154 -3932 1229 -3924
rect 1834 -4026 1896 -3713
rect 2160 -3718 2212 -3712
rect 2326 -3743 2335 -3680
rect 2398 -3743 2780 -3680
rect 2160 -3776 2212 -3770
rect 848 -4033 900 -4027
rect 848 -4091 900 -4085
rect 2717 -3996 2780 -3743
rect 2717 -4065 2780 -4059
rect 1834 -4094 1896 -4088
rect 3375 -4494 3479 -4488
rect 3479 -4598 3559 -4494
rect 3663 -4598 3672 -4494
rect 3375 -4604 3479 -4598
<< via2 >>
rect 627 -3113 687 -3112
rect 627 -3172 686 -3113
rect 686 -3172 687 -3113
rect 1459 -3170 1515 -3114
rect 3228 -3370 3288 -3310
rect 1163 -3921 1219 -3865
rect 2335 -3743 2398 -3680
rect 3559 -4598 3663 -4494
<< metal3 >>
rect 622 -3112 692 -3107
rect 1454 -3112 1520 -3109
rect 622 -3172 627 -3112
rect 687 -3114 1520 -3112
rect 687 -3170 1459 -3114
rect 1515 -3170 1520 -3114
rect 687 -3172 1520 -3170
rect 622 -3177 692 -3172
rect 1454 -3175 1520 -3172
rect 3223 -3310 3293 -3305
rect 3378 -3310 3384 -3308
rect 3223 -3370 3228 -3310
rect 3288 -3370 3384 -3310
rect 3223 -3375 3293 -3370
rect 3378 -3372 3384 -3370
rect 3448 -3372 3454 -3308
rect 2330 -3679 2403 -3675
rect 1159 -3680 2403 -3679
rect 1159 -3742 2335 -3680
rect 1159 -3860 1222 -3742
rect 2330 -3743 2335 -3742
rect 2398 -3743 2403 -3680
rect 2330 -3748 2403 -3743
rect 1158 -3865 1224 -3860
rect 1158 -3921 1163 -3865
rect 1219 -3921 1224 -3865
rect 1158 -3926 1224 -3921
rect 3554 -4494 3668 -4489
rect 3554 -4598 3559 -4494
rect 3663 -4598 3729 -4494
rect 3833 -4598 3839 -4494
rect 3554 -4603 3668 -4598
<< via3 >>
rect 3384 -3372 3448 -3308
rect 3729 -4598 3833 -4494
<< metal4 >>
rect 3383 -3308 3449 -3307
rect 3383 -3372 3384 -3308
rect 3448 -3310 3449 -3308
rect 3448 -3370 3594 -3310
rect 3448 -3372 3449 -3370
rect 3383 -3373 3449 -3372
rect 4185 -4493 4289 -4306
rect 3718 -4494 4289 -4493
rect 3718 -4597 3729 -4494
rect 3728 -4598 3729 -4597
rect 3833 -4597 4289 -4494
rect 3833 -4598 3834 -4597
rect 3728 -4599 3834 -4598
use sky130_fd_pr__cap_mim_m3_1_VLUT89  XC1
timestamp 1755620011
transform 1 0 3900 0 1 -2574
box -386 -1800 386 1800
use sky130_fd_pr__pfet_01v8_XGEKHL  XM1
timestamp 1755620011
transform 1 0 2748 0 1 -3252
box -263 -319 263 319
use sky130_fd_pr__pfet_01v8_XGEKHL  XM6
timestamp 1755620011
transform 1 0 873 0 1 -3250
box -263 -319 263 319
use sky130_fd_pr__nfet_01v8_64Z3AY  XM7
timestamp 1755656603
transform 1 0 821 0 1 -4029
box -211 -279 211 279
use sky130_fd_pr__nfet_01v8_64Z3AY  XM8
timestamp 1755656603
transform 1 0 1812 0 1 -4030
box -211 -279 211 279
use sky130_fd_pr__pfet_01v8_XGEKHL  XM9
timestamp 1755620011
transform 1 0 1867 0 1 -3252
box -263 -319 263 319
use sky130_fd_pr__nfet_01v8_64Z3AY  XM10
timestamp 1755656603
transform 1 0 2801 0 1 -4029
box -211 -279 211 279
<< labels >>
flabel metal2 1834 -4026 1896 -3269 0 FreeSans 320 0 0 0 CLKN
flabel metal2 2717 -3996 2780 -3280 0 FreeSans 320 0 0 0 CLKB
flabel metal1 423 -3740 623 -3540 0 FreeSans 256 0 0 0 SH_IN
port 1 nsew
flabel metal1 424 -4605 624 -4405 0 FreeSans 256 0 0 0 VSS
port 2 nsew
flabel metal1 427 -2830 627 -2630 0 FreeSans 256 0 0 0 VCC
port 3 nsew
flabel metal1 2992 -3737 3192 -3537 0 FreeSans 256 0 0 0 SH_OUT
port 0 nsew
flabel metal1 428 -3243 628 -3043 0 FreeSans 256 0 0 0 SH_CLK
port 4 nsew
<< end >>
