magic
tech sky130A
magscale 1 2
timestamp 1755345873
<< locali >>
rect 7450 -11986 7484 -11852
<< viali >>
rect 6058 -4202 6216 -4168
rect 6734 -4202 6892 -4168
rect 5232 -5142 5266 -5108
rect 4244 -6050 4402 -6016
rect 6060 -6182 6218 -6148
rect 6572 -6182 6730 -6148
rect 5390 -6494 5424 -6460
rect 3410 -6690 3446 -6574
rect 5234 -7116 5268 -7082
rect 6538 -7464 6572 -7378
rect 3502 -7552 3660 -7518
rect 4244 -7548 4402 -7514
rect 5246 -8638 5280 -8604
rect 6918 -8686 7076 -8652
rect 7596 -8684 7754 -8650
rect 6922 -10122 7080 -10088
rect 7500 -10124 7658 -10090
rect 7132 -11868 7170 -11738
<< metal1 >>
rect 6190 -2742 6196 -2740
rect 5684 -2790 6196 -2742
rect 5392 -3844 5452 -3838
rect 5220 -3904 5392 -3844
rect 5220 -4584 5280 -3904
rect 5392 -3910 5452 -3904
rect 4276 -4676 5280 -4584
rect 3527 -5475 3570 -5474
rect 4276 -5475 4368 -4676
rect 5220 -4937 5280 -4676
rect 5554 -4937 5560 -4936
rect 5220 -4987 5560 -4937
rect 5220 -5108 5280 -4987
rect 5554 -4988 5560 -4987
rect 5612 -4988 5618 -4936
rect 5220 -5142 5232 -5108
rect 5266 -5132 5280 -5108
rect 5266 -5142 5278 -5132
rect 5220 -5154 5278 -5142
rect 5212 -5248 5282 -5182
rect 3191 -5518 4368 -5475
rect 3191 -6626 3234 -5518
rect 3527 -5936 3570 -5518
rect 4276 -5582 4368 -5518
rect 4732 -5425 4932 -5334
rect 4732 -5495 5037 -5425
rect 5107 -5495 5227 -5425
rect 4732 -5534 4932 -5495
rect 5279 -5515 5513 -5445
rect 4270 -5674 4276 -5582
rect 4368 -5674 4374 -5582
rect 4770 -5584 4818 -5534
rect 4768 -5590 4820 -5584
rect 4768 -5648 4820 -5642
rect 3915 -5801 3921 -5731
rect 3991 -5801 5287 -5731
rect 4276 -5876 4368 -5870
rect 3360 -6004 4164 -5936
rect 3360 -6376 3428 -6004
rect 3548 -6174 3620 -6106
rect 3921 -6239 3991 -6233
rect 3921 -6373 3991 -6309
rect 3360 -6444 3560 -6376
rect 3607 -6443 3991 -6373
rect 4096 -6370 4164 -6004
rect 4232 -5968 4276 -5924
rect 4368 -5968 4416 -5924
rect 4232 -6016 4416 -5968
rect 4232 -6050 4244 -6016
rect 4402 -6050 4416 -6016
rect 4232 -6062 4416 -6050
rect 4284 -6170 4356 -6102
rect 4668 -6367 4738 -6366
rect 4096 -6438 4306 -6370
rect 4345 -6437 4738 -6367
rect 3388 -6574 3468 -6560
rect 3388 -6626 3410 -6574
rect 3191 -6669 3410 -6626
rect 3388 -6690 3410 -6669
rect 3446 -6690 3468 -6574
rect 3388 -6718 3468 -6690
rect 3548 -6796 3618 -6640
rect 3482 -6996 3682 -6796
rect 3921 -6859 3991 -6443
rect 4290 -6859 4354 -6636
rect 3921 -6929 4354 -6859
rect 3548 -7148 3618 -6996
rect 3921 -7246 3991 -6929
rect 4290 -7142 4354 -6929
rect 4668 -6799 4738 -6437
rect 4903 -6423 4973 -5801
rect 5443 -6050 5513 -5515
rect 5684 -6050 5732 -2790
rect 6190 -2792 6196 -2790
rect 6248 -2792 6254 -2740
rect 6440 -3830 6640 -3764
rect 5942 -3844 6002 -3838
rect 6440 -3844 7703 -3830
rect 6002 -3899 7703 -3844
rect 6002 -3904 6640 -3899
rect 5942 -3910 6002 -3904
rect 6440 -3964 6640 -3904
rect 6440 -4154 6504 -3964
rect 6048 -4168 6910 -4154
rect 6048 -4202 6058 -4168
rect 6216 -4202 6734 -4168
rect 6892 -4202 6910 -4168
rect 6048 -4218 6910 -4202
rect 6104 -4310 6170 -4254
rect 6440 -4612 6504 -4218
rect 6780 -4310 6846 -4254
rect 6158 -4792 6790 -4612
rect 6836 -4794 7202 -4738
rect 6064 -5185 6098 -5013
rect 5955 -5192 6098 -5185
rect 5955 -5194 6188 -5192
rect 5955 -5235 6886 -5194
rect 5955 -5888 6005 -5235
rect 6064 -5250 6886 -5235
rect 6104 -5252 6886 -5250
rect 6106 -5780 6172 -5720
rect 6618 -5776 6684 -5720
rect 7118 -5744 7174 -4794
rect 7010 -5884 7210 -5744
rect 5955 -5938 6114 -5888
rect 6166 -5936 6624 -5888
rect 5443 -6098 6174 -6050
rect 5214 -6186 5284 -6116
rect 5443 -6276 5513 -6098
rect 6036 -6148 6230 -6136
rect 6036 -6182 6060 -6148
rect 6218 -6149 6230 -6148
rect 6272 -6149 6278 -6139
rect 6218 -6182 6278 -6149
rect 6036 -6194 6230 -6182
rect 6272 -6191 6278 -6182
rect 6330 -6191 6336 -6139
rect 6372 -6222 6420 -5936
rect 6674 -5944 7210 -5884
rect 6858 -6038 6918 -5944
rect 6618 -6098 6918 -6038
rect 6630 -6138 6682 -6132
rect 6554 -6148 6630 -6138
rect 6682 -6148 6748 -6138
rect 6554 -6182 6572 -6148
rect 6730 -6182 6748 -6148
rect 6554 -6190 6630 -6182
rect 6682 -6190 6748 -6182
rect 6554 -6196 6748 -6190
rect 5031 -6346 5037 -6276
rect 5107 -6346 5222 -6276
rect 5274 -6346 5513 -6276
rect 6100 -6270 6420 -6222
rect 4903 -6499 4973 -6493
rect 5217 -6799 5287 -6455
rect 5378 -6460 5448 -6448
rect 5378 -6494 5390 -6460
rect 5424 -6494 5448 -6460
rect 5378 -6506 5448 -6494
rect 4668 -6869 5287 -6799
rect 5380 -6812 5436 -6506
rect 3359 -7316 3555 -7249
rect 3604 -7316 3991 -7246
rect 3359 -7662 3426 -7316
rect 4079 -7320 4298 -7250
rect 4668 -7252 4738 -6869
rect 5380 -6874 5436 -6868
rect 6100 -6918 6148 -6270
rect 6364 -6478 6430 -6422
rect 6100 -6966 6372 -6918
rect 5554 -6993 5560 -6992
rect 5230 -7032 5560 -6993
rect 5222 -7043 5560 -7032
rect 5222 -7082 5280 -7043
rect 5554 -7044 5560 -7043
rect 5612 -7044 5618 -6992
rect 5222 -7116 5234 -7082
rect 5268 -7116 5280 -7082
rect 5222 -7128 5280 -7116
rect 4897 -7231 4903 -7161
rect 4973 -7231 5283 -7161
rect 3548 -7466 3614 -7410
rect 3490 -7513 3672 -7506
rect 3852 -7513 3858 -7504
rect 3490 -7518 3858 -7513
rect 3490 -7552 3502 -7518
rect 3660 -7547 3858 -7518
rect 3660 -7552 3672 -7547
rect 3490 -7564 3672 -7552
rect 3852 -7556 3858 -7547
rect 3910 -7556 3916 -7504
rect 4081 -7662 4148 -7320
rect 4346 -7322 4738 -7252
rect 5374 -7274 5380 -7218
rect 5436 -7274 5618 -7218
rect 4290 -7462 4356 -7406
rect 4292 -7502 4344 -7498
rect 4234 -7504 4416 -7502
rect 4234 -7514 4292 -7504
rect 4344 -7514 4416 -7504
rect 4234 -7548 4244 -7514
rect 4402 -7548 4416 -7514
rect 4234 -7556 4292 -7548
rect 4344 -7556 4416 -7548
rect 4234 -7560 4416 -7556
rect 4292 -7562 4344 -7560
rect 3359 -7681 4148 -7662
rect 4301 -7681 4335 -7562
rect 3359 -7715 4335 -7681
rect 3359 -7729 4148 -7715
rect 4301 -13083 4335 -7715
rect 4665 -8153 4735 -7322
rect 4768 -7480 4820 -7474
rect 4983 -7482 5223 -7471
rect 4820 -7530 5223 -7482
rect 5279 -7505 5469 -7435
rect 4768 -7538 4820 -7532
rect 4983 -7541 5223 -7530
rect 4983 -7977 5053 -7541
rect 5216 -7778 5286 -7708
rect 5399 -7977 5469 -7505
rect 5562 -7744 5618 -7274
rect 6420 -7378 6584 -7302
rect 6420 -7388 6538 -7378
rect 6418 -7464 6538 -7388
rect 6572 -7388 6584 -7378
rect 6691 -7388 6733 -6196
rect 6572 -7464 6750 -7388
rect 6418 -7508 6750 -7464
rect 6420 -7520 6584 -7508
rect 5562 -7806 5618 -7800
rect 4977 -8047 4983 -7977
rect 5053 -8047 5059 -7977
rect 5399 -8035 5845 -7977
rect 4665 -8223 5293 -8153
rect 5399 -8322 5469 -8035
rect 5556 -8212 5562 -8156
rect 5618 -8212 5624 -8156
rect 4977 -8400 4983 -8330
rect 5053 -8400 5235 -8330
rect 5288 -8392 5469 -8322
rect 5228 -8568 5298 -8498
rect 5238 -8604 5290 -8598
rect 5182 -8638 5246 -8604
rect 5280 -8638 5340 -8604
rect 5238 -8662 5290 -8638
rect 5238 -8788 5278 -8662
rect 5562 -8788 5618 -8212
rect 5238 -8844 5618 -8788
rect 5787 -8435 5845 -8035
rect 5995 -8435 6053 -8429
rect 5787 -8493 5995 -8435
rect 5238 -13083 5278 -8844
rect 5787 -10174 5845 -8493
rect 5995 -8499 6053 -8493
rect 6169 -10174 6227 -10168
rect 5787 -10232 6169 -10174
rect 6169 -10238 6227 -10232
rect 6364 -10764 6432 -8142
rect 6630 -8770 6750 -7508
rect 7634 -8636 7703 -3899
rect 6906 -8650 7766 -8636
rect 6906 -8652 7596 -8650
rect 6906 -8686 6918 -8652
rect 7076 -8684 7596 -8652
rect 7754 -8684 7766 -8650
rect 7076 -8686 7766 -8684
rect 6906 -8702 7766 -8686
rect 6500 -8890 6750 -8770
rect 6964 -8794 7030 -8738
rect 6500 -10089 6620 -8890
rect 7293 -9094 7359 -8702
rect 7642 -8792 7708 -8736
rect 7022 -9320 7652 -9094
rect 7698 -9320 8096 -9096
rect 6930 -9676 6976 -9634
rect 6930 -9689 7722 -9676
rect 6780 -9728 7722 -9689
rect 6780 -9956 6819 -9728
rect 6930 -9734 7722 -9728
rect 6773 -9962 6825 -9956
rect 6773 -10020 6825 -10014
rect 6910 -10088 7692 -10078
rect 6910 -10089 6922 -10088
rect 6500 -10122 6922 -10089
rect 7080 -10090 7692 -10088
rect 7080 -10122 7500 -10090
rect 6500 -10124 7500 -10122
rect 7658 -10124 7692 -10090
rect 6500 -10130 7692 -10124
rect 6500 -10358 6620 -10130
rect 6910 -10142 7692 -10130
rect 6671 -10232 6677 -10174
rect 6735 -10232 7036 -10174
rect 7546 -10232 7612 -10176
rect 6742 -10448 6748 -10372
rect 6824 -10448 6982 -10372
rect 7026 -10398 7554 -10336
rect 7944 -10340 8096 -9320
rect 6500 -10484 6620 -10478
rect 6968 -10548 7034 -10492
rect 7251 -10663 7313 -10398
rect 7602 -10492 7642 -10434
rect 7944 -10492 8144 -10340
rect 7546 -10540 8144 -10492
rect 7546 -10544 7960 -10540
rect 7251 -10725 7639 -10663
rect 6276 -10854 6476 -10764
rect 6276 -10914 7348 -10854
rect 6276 -10964 6476 -10914
rect 7577 -11147 7639 -10725
rect 7327 -11209 7639 -11147
rect 6494 -11348 6500 -11228
rect 6620 -11348 6626 -11228
rect 6500 -11740 6620 -11348
rect 7042 -11738 7286 -11600
rect 7042 -11740 7132 -11738
rect 6500 -11860 7132 -11740
rect 6500 -13062 6620 -11860
rect 7042 -11868 7132 -11860
rect 7170 -11868 7286 -11738
rect 7042 -12010 7286 -11868
rect 7276 -12630 7342 -12574
rect 9430 -13062 9630 -13006
rect 6500 -13083 9630 -13062
rect 4301 -13090 9630 -13083
rect 9844 -13090 9948 -13084
rect 4301 -13117 9844 -13090
rect 6500 -13182 9844 -13117
rect 9430 -13194 9844 -13182
rect 9430 -13206 9630 -13194
rect 9844 -13200 9948 -13194
<< via1 >>
rect 5392 -3904 5452 -3844
rect 5560 -4988 5612 -4936
rect 5037 -5495 5107 -5425
rect 4276 -5674 4368 -5582
rect 4768 -5642 4820 -5590
rect 3921 -5801 3991 -5731
rect 3921 -6309 3991 -6239
rect 4276 -5968 4368 -5876
rect 6196 -2792 6248 -2740
rect 5942 -3904 6002 -3844
rect 6278 -6191 6330 -6139
rect 6630 -6148 6682 -6138
rect 6630 -6182 6682 -6148
rect 6630 -6190 6682 -6182
rect 5037 -6346 5107 -6276
rect 4903 -6493 4973 -6423
rect 5380 -6868 5436 -6812
rect 5560 -7044 5612 -6992
rect 4903 -7231 4973 -7161
rect 3858 -7556 3910 -7504
rect 5380 -7274 5436 -7218
rect 4292 -7514 4344 -7504
rect 4292 -7548 4344 -7514
rect 4292 -7556 4344 -7548
rect 4768 -7532 4820 -7480
rect 5562 -7800 5618 -7744
rect 4983 -8047 5053 -7977
rect 5562 -8212 5618 -8156
rect 4983 -8400 5053 -8330
rect 5995 -8493 6053 -8435
rect 6169 -10232 6227 -10174
rect 6773 -10014 6825 -9962
rect 6677 -10232 6735 -10174
rect 6500 -10478 6620 -10358
rect 6748 -10448 6824 -10372
rect 6500 -11348 6620 -11228
rect 9844 -13194 9948 -13090
<< metal2 >>
rect 6196 -2740 6248 -2734
rect 6835 -2742 6844 -2736
rect 6248 -2790 6844 -2742
rect 6196 -2798 6248 -2792
rect 6835 -2796 6844 -2790
rect 6904 -2796 6913 -2736
rect 5386 -3904 5392 -3844
rect 5452 -3904 5942 -3844
rect 6002 -3904 6008 -3844
rect 5560 -4936 5612 -4930
rect 5560 -4994 5612 -4988
rect 5037 -5425 5107 -5419
rect 4276 -5582 4368 -5576
rect 4762 -5642 4768 -5590
rect 4820 -5642 4826 -5590
rect 3914 -5731 3998 -5724
rect 3914 -5801 3921 -5731
rect 3991 -5801 3998 -5731
rect 3914 -5802 3998 -5801
rect 3921 -6239 3991 -5802
rect 4276 -5876 4368 -5674
rect 4270 -5968 4276 -5876
rect 4368 -5968 4374 -5876
rect 3915 -6309 3921 -6239
rect 3991 -6309 3997 -6239
rect 4770 -7480 4818 -5642
rect 5037 -6276 5107 -5495
rect 5037 -6352 5107 -6346
rect 4897 -6493 4903 -6423
rect 4973 -6493 4979 -6423
rect 4903 -7161 4973 -6493
rect 5374 -6868 5380 -6812
rect 5436 -6868 5442 -6812
rect 4903 -7237 4973 -7231
rect 5380 -7218 5436 -6868
rect 5561 -6986 5611 -4994
rect 6278 -6139 6330 -6133
rect 6624 -6148 6630 -6138
rect 6330 -6181 6630 -6148
rect 6624 -6190 6630 -6181
rect 6682 -6190 6688 -6138
rect 6278 -6197 6330 -6191
rect 5560 -6992 5612 -6986
rect 5560 -7050 5612 -7044
rect 5380 -7280 5436 -7274
rect 3858 -7504 3910 -7498
rect 4286 -7513 4292 -7504
rect 3910 -7547 4292 -7513
rect 4286 -7556 4292 -7547
rect 4344 -7556 4350 -7504
rect 4762 -7532 4768 -7480
rect 4820 -7532 4826 -7480
rect 3858 -7562 3910 -7556
rect 5556 -7800 5562 -7744
rect 5618 -7800 5624 -7744
rect 4983 -7977 5053 -7971
rect 4983 -8330 5053 -8047
rect 5562 -8156 5618 -7800
rect 5562 -8218 5618 -8212
rect 4983 -8406 5053 -8400
rect 6963 -8435 6972 -8434
rect 5989 -8493 5995 -8435
rect 6053 -8493 6972 -8435
rect 6963 -8494 6972 -8493
rect 7032 -8494 7041 -8434
rect 6767 -10014 6773 -9962
rect 6825 -10014 6831 -9962
rect 6677 -10174 6735 -10168
rect 6163 -10232 6169 -10174
rect 6227 -10232 6677 -10174
rect 6677 -10238 6735 -10232
rect 6494 -10478 6500 -10358
rect 6620 -10478 6626 -10358
rect 6779 -10366 6818 -10014
rect 6748 -10372 6824 -10366
rect 6748 -10454 6824 -10448
rect 6500 -11228 6620 -10478
rect 6500 -11354 6620 -11348
rect 10131 -13090 10225 -13086
rect 9838 -13194 9844 -13090
rect 9948 -13095 10230 -13090
rect 9948 -13189 10131 -13095
rect 10225 -13189 10230 -13095
rect 9948 -13194 10230 -13189
rect 10131 -13198 10225 -13194
<< via2 >>
rect 6844 -2796 6904 -2736
rect 6972 -8494 7032 -8434
rect 10131 -13189 10225 -13095
<< metal3 >>
rect 6839 -2736 6909 -2731
rect 7000 -2736 7006 -2734
rect 6839 -2796 6844 -2736
rect 6904 -2796 7006 -2736
rect 6839 -2801 6909 -2796
rect 7000 -2798 7006 -2796
rect 7070 -2798 7076 -2734
rect 6967 -8434 7037 -8429
rect 7396 -8434 7402 -8432
rect 6967 -8494 6972 -8434
rect 7032 -8494 7402 -8434
rect 6967 -8499 7037 -8494
rect 7396 -8496 7402 -8494
rect 7466 -8496 7472 -8432
rect 10443 -13090 10545 -13085
rect 10126 -13091 10546 -13090
rect 10126 -13095 10443 -13091
rect 10126 -13189 10131 -13095
rect 10225 -13189 10443 -13095
rect 10126 -13193 10443 -13189
rect 10545 -13193 10546 -13091
rect 10126 -13194 10546 -13193
rect 10443 -13199 10545 -13194
<< via3 >>
rect 7006 -2798 7070 -2734
rect 7402 -8496 7466 -8432
rect 10443 -13193 10545 -13091
<< metal4 >>
rect 7005 -2734 7071 -2733
rect 7005 -2798 7006 -2734
rect 7070 -2736 7071 -2734
rect 7070 -2796 8514 -2736
rect 7070 -2798 7071 -2796
rect 7005 -2799 7071 -2798
rect 9062 -5448 9166 -5158
rect 9062 -5552 10548 -5448
rect 10444 -6168 10548 -5552
rect 7404 -8276 9290 -8216
rect 7404 -8431 7464 -8276
rect 7401 -8432 7467 -8431
rect 7401 -8496 7402 -8432
rect 7466 -8496 7467 -8432
rect 7401 -8497 7467 -8496
rect 10442 -13091 10546 -12536
rect 10442 -13193 10443 -13091
rect 10545 -13193 10546 -13091
rect 10442 -13194 10546 -13193
use sky130_fd_pr__pfet_01v8_XGAKDL  sky130_fd_pr__pfet_01v8_XGAKDL_0
timestamp 1755275318
transform 1 0 3585 0 1 -6403
box -211 -419 211 419
use sky130_fd_pr__cap_mim_m3_1_VLUT89  XC1
timestamp 1755275318
transform 1 0 8784 0 1 -3460
box -386 -1800 386 1800
use sky130_fd_pr__cap_mim_m3_1_VLKC9S  XC2
timestamp 1755275318
transform 1 0 9860 0 1 -9246
box -686 -3300 686 3300
use sky130_fd_pr__nfet_01v8_648S5X  XM1
timestamp 1755275318
transform 1 0 6139 0 1 -5908
box -211 -310 211 310
use sky130_fd_pr__nfet_01v8_648S5X  XM2
timestamp 1755275318
transform 1 0 6651 0 1 -5908
box -211 -310 211 310
use sky130_fd_pr__nfet_01v8_QLNS5P  XM3
timestamp 1755275318
transform 1 0 6397 0 1 -7310
box -211 -1010 211 1010
use sky130_fd_pr__pfet_01v8_XGASDL  XM4
timestamp 1755275318
transform 1 0 6137 0 1 -4751
box -211 -619 211 619
use sky130_fd_pr__pfet_01v8_XGASDL  XM5
timestamp 1755275318
transform 1 0 6813 0 1 -4751
box -211 -619 211 619
use sky130_fd_pr__pfet_01v8_XGAKDL  XM6
timestamp 1755275318
transform 1 0 5249 0 1 -5491
box -211 -419 211 419
use sky130_fd_pr__nfet_01v8_648S5X  XM7
timestamp 1755275318
transform 1 0 5249 0 1 -6316
box -211 -310 211 310
use sky130_fd_pr__nfet_01v8_648S5X  XM8
timestamp 1755275318
transform 1 0 3581 0 1 -7278
box -211 -310 211 310
use sky130_fd_pr__nfet_01v8_648S5X  XM10
timestamp 1755275318
transform 1 0 4323 0 1 -7274
box -211 -310 211 310
use sky130_fd_pr__pfet_01v8_XGAKDL  XM11
timestamp 1755275318
transform 1 0 4323 0 1 -6399
box -211 -419 211 419
use sky130_fd_pr__nfet_01v8_648S5X  XM12
timestamp 1755275318
transform 1 0 7001 0 1 -10362
box -211 -310 211 310
use sky130_fd_pr__nfet_01v8_648S5X  XM13
timestamp 1755275318
transform 1 0 7579 0 1 -10364
box -211 -310 211 310
use sky130_fd_pr__nfet_01v8_QLNS5P  XM14
timestamp 1755275318
transform 1 0 7309 0 1 -11742
box -211 -1010 211 1010
use sky130_fd_pr__pfet_01v8_XGASDL  XM15
timestamp 1755275318
transform 1 0 6997 0 1 -9235
box -211 -619 211 619
use sky130_fd_pr__pfet_01v8_XGASDL  XM16
timestamp 1755275318
transform 1 0 7675 0 1 -9233
box -211 -619 211 619
use sky130_fd_pr__pfet_01v8_XGAKDL  XM17
timestamp 1755275318
transform 1 0 5251 0 1 -7465
box -211 -419 211 419
use sky130_fd_pr__nfet_01v8_648S5X  XM18
timestamp 1755275318
transform 1 0 5261 0 1 -8364
box -211 -310 211 310
<< labels >>
flabel metal1 3482 -6996 3682 -6796 0 FreeSans 256 0 0 0 CLK
port 6 nsew
flabel metal1 3921 -6929 4354 -6859 0 FreeSans 800 0 0 0 CLKN
flabel space 4669 -7322 4739 -6367 0 FreeSans 800 0 0 0 CLKB
flabel metal1 4732 -5534 4932 -5334 0 FreeSans 256 0 0 0 SH_IN
port 1 nsew
flabel metal1 7010 -5944 7210 -5744 0 FreeSans 256 0 0 0 SH_OUT
port 0 nsew
flabel metal1 6276 -10964 6476 -10764 0 FreeSans 256 0 0 0 VREF
port 4 nsew
flabel metal1 5787 -10232 5845 -7977 0 FreeSans 800 0 0 0 CIN2
flabel metal1 5684 -6098 5732 -2742 0 FreeSans 800 0 0 0 CIN1
flabel metal1 9430 -13206 9630 -13006 0 FreeSans 256 0 0 0 VSS
port 3 nsew
flabel metal1 6440 -3964 6640 -3764 0 FreeSans 256 0 0 0 VCC
port 5 nsew
flabel metal1 7944 -10540 8144 -10340 0 FreeSans 256 0 0 0 SH_OUT2
port 2 nsew
<< end >>
