magic
tech sky130A
magscale 1 2
timestamp 1761841071
<< metal1 >>
rect 25182 33156 25254 33162
rect 24590 32332 24662 32338
rect 23988 31520 24060 31526
rect 23388 30704 23460 30710
rect 22788 29886 22860 29892
rect 22172 29062 22244 29068
rect 21566 28174 21572 28246
rect 21644 28174 21650 28246
rect 20972 27366 20978 27438
rect 21050 27366 21056 27438
rect 20978 26148 21050 27366
rect 21572 26132 21644 28174
rect 22172 26042 22244 28990
rect 22788 26124 22860 29814
rect 23388 26140 23460 30632
rect 23988 26080 24060 31448
rect 24590 26034 24662 32260
rect 25182 26064 25254 33084
rect 19562 24698 19962 24704
rect 19962 24298 20234 24698
rect 19562 24292 19962 24298
rect 20018 17458 20218 24298
rect 18718 16516 18724 16716
rect 18924 16516 19472 16716
rect 25270 16120 25330 16126
rect 25270 16054 25330 16060
rect 25571 15539 25623 15545
rect 25283 15488 25571 15539
rect 25571 15481 25623 15487
rect 25883 14776 26030 20604
rect 26611 15486 26617 15538
rect 26669 15537 26675 15538
rect 26669 15486 27123 15537
rect 25207 14629 26030 14776
rect 16956 14044 17012 14050
rect 17012 13988 17386 14044
rect 16956 13982 17012 13988
rect 17154 12912 17160 12972
rect 17220 12912 17458 12972
rect 17507 10557 17513 10756
rect 17712 10557 17718 10756
rect 23836 8591 23842 8791
rect 24042 8591 24480 8791
rect 24310 8308 24370 8314
rect 24310 8242 24370 8248
rect 27072 7835 27123 15486
rect 24268 7644 24448 7778
rect 24262 7464 24268 7644
rect 24448 7464 24454 7644
rect 23934 6816 23940 7016
rect 24140 6816 24490 7016
<< via1 >>
rect 25182 33084 25254 33156
rect 24590 32260 24662 32332
rect 23988 31448 24060 31520
rect 23388 30632 23460 30704
rect 22788 29814 22860 29886
rect 22172 28990 22244 29062
rect 21572 28174 21644 28246
rect 20978 27366 21050 27438
rect 19562 24298 19962 24698
rect 18724 16516 18924 16716
rect 25270 16060 25330 16120
rect 25571 15487 25623 15539
rect 26617 15486 26669 15538
rect 16956 13988 17012 14044
rect 17160 12912 17220 12972
rect 17513 10557 17712 10756
rect 23842 8591 24042 8791
rect 24310 8248 24370 8308
rect 24268 7464 24448 7644
rect 23940 6816 24140 7016
<< metal2 >>
rect 5540 42552 5600 42561
rect 5540 42483 5600 42492
rect 5542 41648 5598 42483
rect 10867 41794 10876 41854
rect 10936 41794 10945 41854
rect 10878 41648 10934 41794
rect 16445 41704 16454 41706
rect 16214 41648 16454 41704
rect 16445 41646 16454 41648
rect 16514 41646 16523 41706
rect 24661 33156 24723 33160
rect 24656 33151 25182 33156
rect 24656 33089 24661 33151
rect 24723 33089 25182 33151
rect 24656 33084 25182 33089
rect 25254 33084 25260 33156
rect 24661 33080 24723 33084
rect 23873 32332 23935 32336
rect 23868 32327 24590 32332
rect 23868 32265 23873 32327
rect 23935 32265 24590 32327
rect 23868 32260 24590 32265
rect 24662 32260 24668 32332
rect 23873 32256 23935 32260
rect 23461 31520 23523 31524
rect 23456 31515 23988 31520
rect 23456 31453 23461 31515
rect 23523 31453 23988 31515
rect 23456 31448 23988 31453
rect 24060 31448 24066 31520
rect 23461 31444 23523 31448
rect 22987 30704 23049 30708
rect 22982 30699 23388 30704
rect 22982 30637 22987 30699
rect 23049 30637 23388 30699
rect 22982 30632 23388 30637
rect 23460 30632 23466 30704
rect 22987 30628 23049 30632
rect 22493 29886 22555 29890
rect 22488 29881 22788 29886
rect 22488 29819 22493 29881
rect 22555 29819 22788 29881
rect 22488 29814 22788 29819
rect 22860 29814 22866 29886
rect 22493 29810 22555 29814
rect 21899 29062 21961 29066
rect 21894 29057 22172 29062
rect 21894 28995 21899 29057
rect 21961 28995 22172 29057
rect 21894 28990 22172 28995
rect 22244 28990 22250 29062
rect 21899 28986 21961 28990
rect 21299 28246 21361 28250
rect 21572 28246 21644 28252
rect 21294 28241 21572 28246
rect 21294 28179 21299 28241
rect 21361 28179 21572 28241
rect 21294 28174 21572 28179
rect 21299 28170 21361 28174
rect 21572 28168 21644 28174
rect 20675 27438 20737 27442
rect 20978 27438 21050 27444
rect 20670 27433 20978 27438
rect 20670 27371 20675 27433
rect 20737 27371 20978 27433
rect 20670 27366 20978 27371
rect 20675 27362 20737 27366
rect 20978 27360 21050 27366
rect 10878 14044 10934 25760
rect 19189 24698 19579 24702
rect 19184 24693 19562 24698
rect 19184 24303 19189 24693
rect 19184 24298 19562 24303
rect 19962 24298 19968 24698
rect 19189 24294 19579 24298
rect 18724 16716 18924 16722
rect 18253 16516 18262 16716
rect 18462 16516 18724 16716
rect 18724 16510 18924 16516
rect 25264 16060 25270 16120
rect 25330 16118 25520 16120
rect 25330 16062 25462 16118
rect 25518 16062 25527 16118
rect 25330 16060 25520 16062
rect 25565 15487 25571 15539
rect 25623 15538 25629 15539
rect 26617 15538 26669 15544
rect 25623 15487 26617 15538
rect 26617 15480 26669 15486
rect 10878 13988 16956 14044
rect 17012 13988 17018 14044
rect 17160 13330 17220 13332
rect 17153 13274 17162 13330
rect 17218 13274 17227 13330
rect 17160 12972 17220 13274
rect 17160 12906 17220 12912
rect 17513 10756 17712 10762
rect 17090 10557 17099 10756
rect 17298 10557 17513 10756
rect 17513 10551 17712 10557
rect 23842 8791 24042 8797
rect 23411 8591 23420 8791
rect 23620 8591 23842 8791
rect 23842 8585 24042 8591
rect 24304 8306 24310 8308
rect 24370 8306 24376 8308
rect 24303 8250 24310 8306
rect 24370 8250 24377 8306
rect 24304 8248 24310 8250
rect 24370 8248 24376 8250
rect 24268 7644 24448 7650
rect 24268 7451 24448 7464
rect 24264 7281 24273 7451
rect 24443 7281 24452 7451
rect 24268 7276 24448 7281
rect 23940 7016 24140 7022
rect 23419 6816 23428 7016
rect 23628 6816 23940 7016
rect 23940 6810 24140 6816
<< via2 >>
rect 5540 42492 5600 42552
rect 10876 41794 10936 41854
rect 16454 41646 16514 41706
rect 24661 33089 24723 33151
rect 23873 32265 23935 32327
rect 23461 31453 23523 31515
rect 22987 30637 23049 30699
rect 22493 29819 22555 29881
rect 21899 28995 21961 29057
rect 21299 28179 21361 28241
rect 20675 27371 20737 27433
rect 19189 24303 19562 24693
rect 19562 24303 19579 24693
rect 18262 16516 18462 16716
rect 25462 16062 25518 16118
rect 17162 13274 17218 13330
rect 17099 10557 17298 10756
rect 23420 8591 23620 8791
rect 24312 8250 24368 8306
rect 24273 7281 24443 7451
rect 23428 6816 23628 7016
<< metal3 >>
rect 28206 44406 28212 44470
rect 28276 44406 28282 44470
rect 5538 42760 5602 42766
rect 5538 42690 5602 42696
rect 5540 42557 5600 42690
rect 5535 42552 5605 42557
rect 5535 42492 5540 42552
rect 5600 42492 5605 42552
rect 5535 42487 5605 42492
rect 10871 41854 10941 41859
rect 28214 41854 28274 44406
rect 28758 44401 28764 44465
rect 28828 44401 28834 44465
rect 10871 41794 10876 41854
rect 10936 41794 28274 41854
rect 10871 41789 10941 41794
rect 16449 41706 16519 41711
rect 28766 41706 28826 44401
rect 16449 41646 16454 41706
rect 16514 41646 28826 41706
rect 16449 41641 16519 41646
rect 18828 39584 19000 39704
rect 19120 39584 19126 39704
rect 18828 38768 19208 38888
rect 19328 38768 19334 38888
rect 18828 37952 19396 38072
rect 19516 37952 19522 38072
rect 18828 37136 19598 37256
rect 19718 37136 19724 37256
rect 18828 36320 19814 36440
rect 19934 36320 19940 36440
rect 18828 35504 20064 35624
rect 20184 35504 20190 35624
rect 18828 34688 20314 34808
rect 20434 34688 20440 34808
rect 18828 33872 20572 33992
rect 20692 33872 20698 33992
rect 18886 33151 24728 33156
rect 18886 33089 24661 33151
rect 24723 33089 24728 33151
rect 18886 33084 24728 33089
rect 18844 32327 23940 32332
rect 18844 32265 23873 32327
rect 23935 32265 23940 32327
rect 18844 32260 23940 32265
rect 18812 31515 23528 31520
rect 18812 31453 23461 31515
rect 23523 31453 23528 31515
rect 18812 31448 23528 31453
rect 18870 30699 23054 30704
rect 18870 30637 22987 30699
rect 23049 30637 23054 30699
rect 18870 30632 23054 30637
rect 18828 29881 22560 29886
rect 18828 29819 22493 29881
rect 22555 29819 22560 29881
rect 18828 29814 22560 29819
rect 18844 29057 21966 29062
rect 18844 28995 21899 29057
rect 21961 28995 21966 29057
rect 18844 28990 21966 28995
rect 18752 28241 21366 28246
rect 18752 28179 21299 28241
rect 21361 28179 21366 28241
rect 18752 28174 21366 28179
rect 18828 27433 20742 27438
rect 18828 27371 20675 27433
rect 20737 27371 20742 27433
rect 18828 27366 20742 27371
rect 5173 25435 5528 25441
rect 8885 25435 9240 25441
rect 222 25431 5171 25435
rect 219 25081 225 25431
rect 575 25081 5171 25431
rect 222 25078 5171 25081
rect 5528 25078 8883 25435
rect 9240 25078 12575 25435
rect 12932 25078 16273 25435
rect 16630 25078 16636 25435
rect 5173 25072 5528 25078
rect 8885 25072 9240 25078
rect 18639 24698 19037 24703
rect 18638 24697 19584 24698
rect 18638 24299 18639 24697
rect 19037 24693 19584 24697
rect 19037 24303 19189 24693
rect 19579 24303 19584 24693
rect 19037 24299 19584 24303
rect 18638 24298 19584 24299
rect 18639 24293 19037 24298
rect 17158 17060 17222 17066
rect 17158 16990 17222 16996
rect 17160 13335 17220 16990
rect 18257 16716 18467 16721
rect 17960 16516 17966 16716
rect 18166 16516 18262 16716
rect 18462 16516 18467 16716
rect 18257 16511 18467 16516
rect 25457 16120 25523 16123
rect 25670 16122 25734 16128
rect 25457 16118 25670 16120
rect 25457 16062 25462 16118
rect 25518 16062 25670 16118
rect 25457 16060 25670 16062
rect 25457 16057 25523 16060
rect 25670 16052 25734 16058
rect 17157 13330 17223 13335
rect 17157 13274 17162 13330
rect 17218 13274 17223 13330
rect 17157 13269 17223 13274
rect 28766 11006 28826 41646
rect 26136 10946 28826 11006
rect 17094 10756 17303 10761
rect 315 10557 321 10756
rect 520 10557 17099 10756
rect 17298 10557 17303 10756
rect 17094 10552 17303 10557
rect 26136 9628 26196 10946
rect 24310 9568 26196 9628
rect 23415 8791 23625 8796
rect 308 8591 314 8791
rect 514 8591 23420 8791
rect 23620 8591 23625 8791
rect 23415 8586 23625 8591
rect 24310 8311 24370 9568
rect 24307 8306 24373 8311
rect 24307 8250 24312 8306
rect 24368 8250 24373 8306
rect 24307 8245 24373 8250
rect 24268 7451 24448 7456
rect 24268 7281 24273 7451
rect 24443 7281 24448 7451
rect 24268 7239 24448 7281
rect 24268 7061 24269 7239
rect 24447 7061 24448 7239
rect 24268 7060 24448 7061
rect 24269 7055 24447 7060
rect 23423 7016 23633 7021
rect 22838 6816 22844 7016
rect 23044 6816 23428 7016
rect 23628 6816 23633 7016
rect 23423 6811 23633 6816
rect 378 2815 384 3015
rect 584 2815 1818 3015
<< via3 >>
rect 28212 44406 28276 44470
rect 5538 42696 5602 42760
rect 28764 44401 28828 44465
rect 19000 39584 19120 39704
rect 19208 38768 19328 38888
rect 19396 37952 19516 38072
rect 19598 37136 19718 37256
rect 19814 36320 19934 36440
rect 20064 35504 20184 35624
rect 20314 34688 20434 34808
rect 20572 33872 20692 33992
rect 225 25081 575 25431
rect 5171 25078 5528 25435
rect 8883 25078 9240 25435
rect 12575 25078 12932 25435
rect 16273 25078 16630 25435
rect 18639 24299 19037 24697
rect 17158 16996 17222 17060
rect 17966 16516 18166 16716
rect 25670 16058 25734 16122
rect 321 10557 520 10756
rect 314 8591 514 8791
rect 24269 7061 24447 7239
rect 22844 6816 23044 7016
rect 384 2815 584 3015
<< metal4 >>
rect 6134 44152 6194 45152
rect 6686 44152 6746 45152
rect 7238 44152 7298 45152
rect 7790 44152 7850 45152
rect 8342 44152 8402 45152
rect 8894 44152 8954 45152
rect 9446 44152 9506 45152
rect 9998 44152 10058 45152
rect 10550 44152 10610 45152
rect 11102 44152 11162 45152
rect 11654 44152 11714 45152
rect 12206 44152 12266 45152
rect 12758 44152 12818 45152
rect 13310 44152 13370 45152
rect 13862 44152 13922 45152
rect 200 25431 600 44152
rect 200 25081 225 25431
rect 575 25081 600 25431
rect 200 10756 600 25081
rect 200 10557 321 10756
rect 520 10557 600 10756
rect 200 8791 600 10557
rect 200 8591 314 8791
rect 514 8591 600 8791
rect 200 3015 600 8591
rect 200 2815 384 3015
rect 584 2815 600 3015
rect 200 1000 600 2815
rect 800 43752 13968 44152
rect 800 24698 1200 43752
rect 14414 43498 14474 45152
rect 5540 43438 14474 43498
rect 5540 42761 5600 43438
rect 5537 42760 5603 42761
rect 5537 42696 5538 42760
rect 5602 42696 5603 42760
rect 5537 42695 5603 42696
rect 14966 42120 15026 45152
rect 15518 42336 15578 45152
rect 16070 42540 16130 45152
rect 16622 42766 16682 45152
rect 17174 42960 17234 45152
rect 17726 43186 17786 45152
rect 18278 43402 18338 45152
rect 18830 43616 18890 45152
rect 19382 44952 19442 45152
rect 19934 44952 19994 45152
rect 20486 44952 20546 45152
rect 21038 44952 21098 45152
rect 21590 44952 21650 45152
rect 22142 44952 22202 45152
rect 22694 44952 22754 45152
rect 23246 44952 23306 45152
rect 23798 44952 23858 45152
rect 24350 44952 24410 45152
rect 24902 44952 24962 45152
rect 25454 44952 25514 45152
rect 26006 44952 26066 45152
rect 26558 44952 26618 45152
rect 18830 43496 20692 43616
rect 18278 43282 20434 43402
rect 17726 43066 20184 43186
rect 17174 42840 19934 42960
rect 16622 42646 19718 42766
rect 16070 42420 19516 42540
rect 15518 42216 19328 42336
rect 14966 42000 19120 42120
rect 19000 39705 19120 42000
rect 18999 39704 19121 39705
rect 18999 39584 19000 39704
rect 19120 39584 19121 39704
rect 18999 39583 19121 39584
rect 19208 38889 19328 42216
rect 19207 38888 19329 38889
rect 19207 38768 19208 38888
rect 19328 38768 19329 38888
rect 19207 38767 19329 38768
rect 19396 38073 19516 42420
rect 19395 38072 19517 38073
rect 19395 37952 19396 38072
rect 19516 37952 19517 38072
rect 19395 37951 19517 37952
rect 19598 37257 19718 42646
rect 19597 37256 19719 37257
rect 19597 37136 19598 37256
rect 19718 37136 19719 37256
rect 19597 37135 19719 37136
rect 19814 36441 19934 42840
rect 19813 36440 19935 36441
rect 19813 36320 19814 36440
rect 19934 36320 19935 36440
rect 19813 36319 19935 36320
rect 20064 35625 20184 43066
rect 20063 35624 20185 35625
rect 20063 35504 20064 35624
rect 20184 35504 20185 35624
rect 20063 35503 20185 35504
rect 20314 34809 20434 43282
rect 20313 34808 20435 34809
rect 20313 34688 20314 34808
rect 20434 34688 20435 34808
rect 20313 34687 20435 34688
rect 20572 33993 20692 43496
rect 20571 33992 20693 33993
rect 20571 33872 20572 33992
rect 20692 33872 20693 33992
rect 20571 33871 20693 33872
rect 5191 25436 5511 26618
rect 5170 25435 5529 25436
rect 5170 25078 5171 25435
rect 5528 25078 5529 25435
rect 5170 25077 5529 25078
rect 7042 24698 7362 26600
rect 8893 25436 9213 26616
rect 8882 25435 9241 25436
rect 8882 25078 8883 25435
rect 9240 25078 9241 25435
rect 8882 25077 9241 25078
rect 10744 24698 11064 26636
rect 12595 25436 12915 26648
rect 12574 25435 12933 25436
rect 12574 25078 12575 25435
rect 12932 25078 12933 25435
rect 12574 25077 12933 25078
rect 14446 24698 14766 26600
rect 16297 25436 16617 26596
rect 16272 25435 16631 25436
rect 16272 25078 16273 25435
rect 16630 25078 16631 25435
rect 16272 25077 16631 25078
rect 800 24697 19038 24698
rect 800 24299 18639 24697
rect 19037 24299 19038 24697
rect 800 24298 19038 24299
rect 800 16716 1200 24298
rect 17157 17060 17223 17061
rect 17157 16996 17158 17060
rect 17222 17058 17223 17060
rect 27110 17058 27170 45152
rect 17222 16998 27170 17058
rect 17222 16996 17223 16998
rect 17157 16995 17223 16996
rect 17965 16716 18167 16717
rect 800 16516 17966 16716
rect 18166 16516 18167 16716
rect 800 7016 1200 16516
rect 17965 16515 18167 16516
rect 25669 16122 25735 16123
rect 25669 16058 25670 16122
rect 25734 16120 25735 16122
rect 27662 16120 27722 45152
rect 28214 44471 28274 45152
rect 28211 44470 28277 44471
rect 28211 44406 28212 44470
rect 28276 44406 28277 44470
rect 28766 44466 28826 45152
rect 29318 44952 29378 45152
rect 28211 44405 28277 44406
rect 28763 44465 28829 44466
rect 28763 44401 28764 44465
rect 28828 44401 28829 44465
rect 28763 44400 28829 44401
rect 25734 16060 27722 16120
rect 25734 16058 25735 16060
rect 25669 16057 25735 16058
rect 24268 7239 24448 7240
rect 24268 7061 24269 7239
rect 24447 7061 24448 7239
rect 22843 7016 23045 7017
rect 800 6816 22844 7016
rect 23044 6816 23045 7016
rect 800 1433 1200 6816
rect 22843 6815 23045 6816
rect 24268 4832 24448 7061
rect 24268 4652 30542 4832
rect 800 1033 1788 1433
rect 800 1000 1200 1033
rect 3314 0 3494 200
rect 7178 0 7358 200
rect 11042 0 11222 200
rect 14906 0 15086 200
rect 18770 0 18950 200
rect 22634 0 22814 200
rect 26498 0 26678 200
rect 30362 0 30542 4652
use comparator  comparator_0
timestamp 1757527180
transform -1 0 31305 0 -1 9227
box 5945 -7489 14005 -1329
use r2r_dac  r2r_dac_0
timestamp 1755981703
transform 1 0 21018 0 1 21522
box -1000 -4230 5038 4682
use Sample_and_Hold  Sample_and_Hold_0
timestamp 1755657154
transform 1 0 23841 0 1 11421
box 423 -4605 4289 -774
use sar_control  sar_control_0
timestamp 1761224974
transform 1 0 2948 0 1 25704
box 514 0 16000 16000
<< labels >>
flabel metal4 s 28766 44952 28826 45152 0 FreeSans 480 90 0 0 clk
port 0 nsew signal input
flabel metal4 s 29318 44952 29378 45152 0 FreeSans 480 90 0 0 ena
port 1 nsew signal input
flabel metal4 s 28214 44952 28274 45152 0 FreeSans 480 90 0 0 rst_n
port 2 nsew signal input
flabel metal4 s 30362 0 30542 200 0 FreeSans 960 0 0 0 ua[0]
port 3 nsew signal bidirectional
flabel metal4 s 26498 0 26678 200 0 FreeSans 960 0 0 0 ua[1]
port 4 nsew signal bidirectional
flabel metal4 s 22634 0 22814 200 0 FreeSans 960 0 0 0 ua[2]
port 5 nsew signal bidirectional
flabel metal4 s 18770 0 18950 200 0 FreeSans 960 0 0 0 ua[3]
port 6 nsew signal bidirectional
flabel metal4 s 14906 0 15086 200 0 FreeSans 960 0 0 0 ua[4]
port 7 nsew signal bidirectional
flabel metal4 s 11042 0 11222 200 0 FreeSans 960 0 0 0 ua[5]
port 8 nsew signal bidirectional
flabel metal4 s 7178 0 7358 200 0 FreeSans 960 0 0 0 ua[6]
port 9 nsew signal bidirectional
flabel metal4 s 3314 0 3494 200 0 FreeSans 960 0 0 0 ua[7]
port 10 nsew signal bidirectional
flabel metal4 s 27662 44952 27722 45152 0 FreeSans 480 90 0 0 ui_in[0]
port 11 nsew signal input
flabel metal4 s 27110 44952 27170 45152 0 FreeSans 480 90 0 0 ui_in[1]
port 12 nsew signal input
flabel metal4 s 26558 44952 26618 45152 0 FreeSans 480 90 0 0 ui_in[2]
port 13 nsew signal input
flabel metal4 s 26006 44952 26066 45152 0 FreeSans 480 90 0 0 ui_in[3]
port 14 nsew signal input
flabel metal4 s 25454 44952 25514 45152 0 FreeSans 480 90 0 0 ui_in[4]
port 15 nsew signal input
flabel metal4 s 24902 44952 24962 45152 0 FreeSans 480 90 0 0 ui_in[5]
port 16 nsew signal input
flabel metal4 s 24350 44952 24410 45152 0 FreeSans 480 90 0 0 ui_in[6]
port 17 nsew signal input
flabel metal4 s 23798 44952 23858 45152 0 FreeSans 480 90 0 0 ui_in[7]
port 18 nsew signal input
flabel metal4 s 23246 44952 23306 45152 0 FreeSans 480 90 0 0 uio_in[0]
port 19 nsew signal input
flabel metal4 s 22694 44952 22754 45152 0 FreeSans 480 90 0 0 uio_in[1]
port 20 nsew signal input
flabel metal4 s 22142 44952 22202 45152 0 FreeSans 480 90 0 0 uio_in[2]
port 21 nsew signal input
flabel metal4 s 21590 44952 21650 45152 0 FreeSans 480 90 0 0 uio_in[3]
port 22 nsew signal input
flabel metal4 s 21038 44952 21098 45152 0 FreeSans 480 90 0 0 uio_in[4]
port 23 nsew signal input
flabel metal4 s 20486 44952 20546 45152 0 FreeSans 480 90 0 0 uio_in[5]
port 24 nsew signal input
flabel metal4 s 19934 44952 19994 45152 0 FreeSans 480 90 0 0 uio_in[6]
port 25 nsew signal input
flabel metal4 s 19382 44952 19442 45152 0 FreeSans 480 90 0 0 uio_in[7]
port 26 nsew signal input
flabel metal4 s 9998 44952 10058 45152 0 FreeSans 480 90 0 0 uio_oe[0]
port 27 nsew signal output
flabel metal4 s 9446 44952 9506 45152 0 FreeSans 480 90 0 0 uio_oe[1]
port 28 nsew signal output
flabel metal4 s 8894 44952 8954 45152 0 FreeSans 480 90 0 0 uio_oe[2]
port 29 nsew signal output
flabel metal4 s 8342 44952 8402 45152 0 FreeSans 480 90 0 0 uio_oe[3]
port 30 nsew signal output
flabel metal4 s 7790 44952 7850 45152 0 FreeSans 480 90 0 0 uio_oe[4]
port 31 nsew signal output
flabel metal4 s 7238 44952 7298 45152 0 FreeSans 480 90 0 0 uio_oe[5]
port 32 nsew signal output
flabel metal4 s 6686 44952 6746 45152 0 FreeSans 480 90 0 0 uio_oe[6]
port 33 nsew signal output
flabel metal4 s 6134 44952 6194 45152 0 FreeSans 480 90 0 0 uio_oe[7]
port 34 nsew signal output
flabel metal4 s 14414 44952 14474 45152 0 FreeSans 480 90 0 0 uio_out[0]
port 35 nsew signal output
flabel metal4 s 13862 44952 13922 45152 0 FreeSans 480 90 0 0 uio_out[1]
port 36 nsew signal output
flabel metal4 s 13310 44952 13370 45152 0 FreeSans 480 90 0 0 uio_out[2]
port 37 nsew signal output
flabel metal4 s 12758 44952 12818 45152 0 FreeSans 480 90 0 0 uio_out[3]
port 38 nsew signal output
flabel metal4 s 12206 44952 12266 45152 0 FreeSans 480 90 0 0 uio_out[4]
port 39 nsew signal output
flabel metal4 s 11654 44952 11714 45152 0 FreeSans 480 90 0 0 uio_out[5]
port 40 nsew signal output
flabel metal4 s 11102 44952 11162 45152 0 FreeSans 480 90 0 0 uio_out[6]
port 41 nsew signal output
flabel metal4 s 10550 44952 10610 45152 0 FreeSans 480 90 0 0 uio_out[7]
port 42 nsew signal output
flabel metal4 s 18830 44952 18890 45152 0 FreeSans 480 90 0 0 uo_out[0]
port 43 nsew signal output
flabel metal4 s 18278 44952 18338 45152 0 FreeSans 480 90 0 0 uo_out[1]
port 44 nsew signal output
flabel metal4 s 17726 44952 17786 45152 0 FreeSans 480 90 0 0 uo_out[2]
port 45 nsew signal output
flabel metal4 s 17174 44952 17234 45152 0 FreeSans 480 90 0 0 uo_out[3]
port 46 nsew signal output
flabel metal4 s 16622 44952 16682 45152 0 FreeSans 480 90 0 0 uo_out[4]
port 47 nsew signal output
flabel metal4 s 16070 44952 16130 45152 0 FreeSans 480 90 0 0 uo_out[5]
port 48 nsew signal output
flabel metal4 s 15518 44952 15578 45152 0 FreeSans 480 90 0 0 uo_out[6]
port 49 nsew signal output
flabel metal4 s 14966 44952 15026 45152 0 FreeSans 480 90 0 0 uo_out[7]
port 50 nsew signal output
flabel metal4 200 1000 600 44152 1 FreeSans 1600 0 0 0 VDPWR
port 51 nsew power bidirectional
flabel metal4 800 1000 1200 44152 1 FreeSans 1600 0 0 0 VGND
port 52 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 32200 45152
<< end >>
