** sch_path: /home/ttuser/ttsky_SAR_ADC/xschem/Sample_and_Hold.sch
.subckt Sample_and_Hold SH_OUT SH_IN VSS VCC SH_CLK
*.PININFO SH_IN:I SH_CLK:I SH_OUT:O VSS:I VCC:I
XC1 SH_OUT VSS sky130_fd_pr__cap_mim_m3_1 W=2 L=2 m=5
XM6 SH_OUT CLKN SH_IN VCC sky130_fd_pr__pfet_01v8 L=0.15 W=2 nf=2 m=1
XM7 SH_IN CLKB SH_OUT VSS sky130_fd_pr__nfet_01v8 L=0.15 W=1 nf=1 m=1
XM8 CLKN SH_CLK VSS VSS sky130_fd_pr__nfet_01v8 L=0.15 W=1 nf=1 m=1
XM9 CLKN SH_CLK VCC VCC sky130_fd_pr__pfet_01v8 L=0.15 W=2 nf=2 m=1
XM10 CLKB CLKN VSS VSS sky130_fd_pr__nfet_01v8 L=0.15 W=1 nf=1 m=1
XM1 CLKB CLKN VCC VCC sky130_fd_pr__pfet_01v8 L=0.15 W=2 nf=2 m=1
.ends
.end
