** sch_path: /home/ttuser/ttsky_SAR_ADC/xschem/Sample_and_Hold.sch
.subckt Sample_and_Hold SH_OUT SH_IN SH_OUT2 VSS VREF VCC CLK
*.PININFO SH_IN:I CLK:I SH_OUT:O VSS:I VCC:I SH_OUT2:O VREF:I
XM1 net2 CIN net1 VSS sky130_fd_pr__nfet_01v8 L=0.15 W=1 nf=1 m=1
XM2 SH_OUT SH_OUT net1 VSS sky130_fd_pr__nfet_01v8 L=0.15 W=1 nf=1 m=1
XM3 net1 VREF VSS VSS sky130_fd_pr__nfet_01v8 L=0.15 W=8 nf=1 m=1
XM4 net2 net2 VCC VCC sky130_fd_pr__pfet_01v8 L=0.15 W=4 nf=1 m=1
XM5 SH_OUT net2 VCC VCC sky130_fd_pr__pfet_01v8 L=0.15 W=4 nf=1 m=1
XC1 CIN VSS sky130_fd_pr__cap_mim_m3_1 W=2 L=2 m=5
XM6 CIN CLKN SH_IN VCC sky130_fd_pr__pfet_01v8 L=0.15 W=2 nf=1 m=1
XM7 SH_IN CLKB CIN VSS sky130_fd_pr__nfet_01v8 L=0.15 W=1 nf=1 m=1
XM8 CLKN CLK VSS VSS sky130_fd_pr__nfet_01v8 L=0.15 W=1 nf=1 m=1
XM9 CLKN CLK VCC VCC sky130_fd_pr__pfet_01v8 L=0.15 W=2 nf=1 m=1
XM10 CLKB CLKN VSS VSS sky130_fd_pr__nfet_01v8 L=0.15 W=1 nf=1 m=1
XM11 CLKB CLKN VCC VCC sky130_fd_pr__pfet_01v8 L=0.15 W=2 nf=1 m=1
XC2 CIN2 VSS sky130_fd_pr__cap_mim_m3_1 W=5 L=5 m=5
XM17 CIN2 CLKN SH_IN VCC sky130_fd_pr__pfet_01v8 L=0.15 W=2 nf=1 m=1
XM18 SH_IN CLKB CIN2 VSS sky130_fd_pr__nfet_01v8 L=0.15 W=1 nf=1 m=1
XM12 net4 CIN2 net3 VSS sky130_fd_pr__nfet_01v8 L=0.15 W=1 nf=1 m=1
XM13 SH_OUT2 SH_OUT2 net3 VSS sky130_fd_pr__nfet_01v8 L=0.15 W=1 nf=1 m=1
XM14 net3 VREF VSS VSS sky130_fd_pr__nfet_01v8 L=0.15 W=8 nf=1 m=1
XM15 net4 net4 VCC VCC sky130_fd_pr__pfet_01v8 L=0.15 W=4 nf=1 m=1
XM16 SH_OUT2 net4 VCC VCC sky130_fd_pr__pfet_01v8 L=0.15 W=4 nf=1 m=1
.ends
.end
