magic
tech sky130A
timestamp 1757456334
<< pwell >>
rect -198 -205 198 205
<< nmoslvt >>
rect -100 -100 100 100
<< ndiff >>
rect -129 94 -100 100
rect -129 -94 -123 94
rect -106 -94 -100 94
rect -129 -100 -100 -94
rect 100 94 129 100
rect 100 -94 106 94
rect 123 -94 129 94
rect 100 -100 129 -94
<< ndiffc >>
rect -123 -94 -106 94
rect 106 -94 123 94
<< psubdiff >>
rect -180 170 -132 187
rect 132 170 180 187
rect -180 139 -163 170
rect 163 139 180 170
rect -180 -170 -163 -139
rect 163 -170 180 -139
rect -180 -187 -132 -170
rect 132 -187 180 -170
<< psubdiffcont >>
rect -132 170 132 187
rect -180 -139 -163 139
rect 163 -139 180 139
rect -132 -187 132 -170
<< poly >>
rect -100 136 100 144
rect -100 119 -92 136
rect 92 119 100 136
rect -100 100 100 119
rect -100 -119 100 -100
rect -100 -136 -92 -119
rect 92 -136 100 -119
rect -100 -144 100 -136
<< polycont >>
rect -92 119 92 136
rect -92 -136 92 -119
<< locali >>
rect -180 170 -132 187
rect 132 170 180 187
rect -180 139 -163 170
rect 163 139 180 170
rect -100 119 -92 136
rect 92 119 100 136
rect -123 94 -106 102
rect -123 -102 -106 -94
rect 106 94 123 102
rect 106 -102 123 -94
rect -100 -136 -92 -119
rect 92 -136 100 -119
rect -180 -170 -163 -139
rect 163 -170 180 -139
rect -180 -187 -132 -170
rect 132 -187 180 -170
<< viali >>
rect -92 119 92 136
rect -123 -94 -106 94
rect 106 -94 123 94
rect -92 -136 92 -119
<< metal1 >>
rect -98 136 98 139
rect -98 119 -92 136
rect 92 119 98 136
rect -98 116 98 119
rect -126 94 -103 100
rect -126 -94 -123 94
rect -106 -94 -103 94
rect -126 -100 -103 -94
rect 103 94 126 100
rect 103 -94 106 94
rect 123 -94 126 94
rect 103 -100 126 -94
rect -98 -119 98 -116
rect -98 -136 -92 -119
rect 92 -136 98 -119
rect -98 -139 98 -136
<< properties >>
string FIXED_BBOX -171 -178 171 178
string gencell sky130_fd_pr__nfet_01v8_lvt
string library sky130
string parameters w 2.0 l 2.0 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
