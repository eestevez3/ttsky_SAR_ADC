/*
 * Copyright (c) 2024 Your Name
 * SPDX-License-Identifier: Apache-2.0
 */

`default_nettype none

module tt_um_eestevez3_SAR_ADC (
    input  wire       VGND,
    input  wire       VDPWR,    // 1.8v power supply
//    input  wire       VAPWR,    // 3.3v power supply
    input  wire [7:0] ui_in,    // Dedicated inputs
    output wire [7:0] uo_out,   // Dedicated outputs
    input  wire [7:0] uio_in,   // IOs: Input path
    output wire [7:0] uio_out,  // IOs: Output path
    output wire [7:0] uio_oe,   // IOs: Enable path (active high: 0=input, 1=output)
    inout  wire [7:0] ua,       // Analog pins, only ua[5:0] can be used
    input  wire       ena,      // always 1 when the design is powered, so you can ignore it
    input  wire       clk,      // clock
    input  wire       rst_n     // reset_n - low to reset
);

	Sample_and_Hold Sample_and_Hold(
		.VCC(VDPWR)
		.VSS(VGND)
		.SH_IN(ua[1])
		.SH_OUT(ua[0])
		.SH_CLK(clk)
	);
	
	comparator comparator(
		.VCC(VDPWR)
		.VSS(VGND)
		.CAL(clk)
		.EN_N(clk)
		.PLUS(ua[2])
		.MINUS(ua[3])
		.COMP_OUT(ua[4])
	);
	
	r2r_dac r2r_dac(
		.VSS(VGND)
		.VSUBS(VGND)
		.b0(ui_in[0])
		.b1(ui_in[1])
		.b2(ui_in[2])
		.b3(ui_in[3])
		.b4(ui_in[4])
		.b5(ui_in[5])
		.b6(ui_in[6])
		.b7(ui_in[7])
		.dac_out([ua[5])
	);
    
    assign uo_out[0] = VGND;
    assign uo_out[1] = VGND;
    assign uo_out[2] = VGND;
    assign uo_out[3] = VGND;
    assign uo_out[4] = VGND;
    assign uo_out[5] = VGND;
    assign uo_out[6] = VGND;
    assign uo_out[7] = VGND;

    assign uio_out[0] = VGND;
    assign uio_out[1] = VGND;
    assign uio_out[2] = VGND;
    assign uio_out[3] = VGND;
    assign uio_out[4] = VGND;
    assign uio_out[5] = VGND;
    assign uio_out[6] = VGND;
    assign uio_out[7] = VGND;

    assign uio_oe[0] = VGND;
    assign uio_oe[1] = VGND;
    assign uio_oe[2] = VGND;
    assign uio_oe[3] = VGND;
    assign uio_oe[4] = VGND;
    assign uio_oe[5] = VGND;
    assign uio_oe[6] = VGND;
    assign uio_oe[7] = VGND;

endmodule
