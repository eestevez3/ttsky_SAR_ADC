magic
tech sky130A
magscale 1 2
timestamp 1755275318
<< metal3 >>
rect -686 3152 686 3180
rect -686 2128 602 3152
rect 666 2128 686 3152
rect -686 2100 686 2128
rect -686 1832 686 1860
rect -686 808 602 1832
rect 666 808 686 1832
rect -686 780 686 808
rect -686 512 686 540
rect -686 -512 602 512
rect 666 -512 686 512
rect -686 -540 686 -512
rect -686 -808 686 -780
rect -686 -1832 602 -808
rect 666 -1832 686 -808
rect -686 -1860 686 -1832
rect -686 -2128 686 -2100
rect -686 -3152 602 -2128
rect 666 -3152 686 -2128
rect -686 -3180 686 -3152
<< via3 >>
rect 602 2128 666 3152
rect 602 808 666 1832
rect 602 -512 666 512
rect 602 -1832 666 -808
rect 602 -3152 666 -2128
<< mimcap >>
rect -646 3100 354 3140
rect -646 2180 -606 3100
rect 314 2180 354 3100
rect -646 2140 354 2180
rect -646 1780 354 1820
rect -646 860 -606 1780
rect 314 860 354 1780
rect -646 820 354 860
rect -646 460 354 500
rect -646 -460 -606 460
rect 314 -460 354 460
rect -646 -500 354 -460
rect -646 -860 354 -820
rect -646 -1780 -606 -860
rect 314 -1780 354 -860
rect -646 -1820 354 -1780
rect -646 -2180 354 -2140
rect -646 -3100 -606 -2180
rect 314 -3100 354 -2180
rect -646 -3140 354 -3100
<< mimcapcontact >>
rect -606 2180 314 3100
rect -606 860 314 1780
rect -606 -460 314 460
rect -606 -1780 314 -860
rect -606 -3100 314 -2180
<< metal4 >>
rect -198 3101 -94 3300
rect 582 3152 686 3300
rect -607 3100 315 3101
rect -607 2180 -606 3100
rect 314 2180 315 3100
rect -607 2179 315 2180
rect -198 1781 -94 2179
rect 582 2128 602 3152
rect 666 2128 686 3152
rect 582 1832 686 2128
rect -607 1780 315 1781
rect -607 860 -606 1780
rect 314 860 315 1780
rect -607 859 315 860
rect -198 461 -94 859
rect 582 808 602 1832
rect 666 808 686 1832
rect 582 512 686 808
rect -607 460 315 461
rect -607 -460 -606 460
rect 314 -460 315 460
rect -607 -461 315 -460
rect -198 -859 -94 -461
rect 582 -512 602 512
rect 666 -512 686 512
rect 582 -808 686 -512
rect -607 -860 315 -859
rect -607 -1780 -606 -860
rect 314 -1780 315 -860
rect -607 -1781 315 -1780
rect -198 -2179 -94 -1781
rect 582 -1832 602 -808
rect 666 -1832 686 -808
rect 582 -2128 686 -1832
rect -607 -2180 315 -2179
rect -607 -3100 -606 -2180
rect 314 -3100 315 -2180
rect -607 -3101 315 -3100
rect -198 -3300 -94 -3101
rect 582 -3152 602 -2128
rect 666 -3152 686 -2128
rect 582 -3300 686 -3152
<< properties >>
string FIXED_BBOX -686 2100 394 3180
string gencell sky130_fd_pr__cap_mim_m3_1
string library sky130
string parameters w 5.0 l 5.0 val 53.8 carea 2.00 cperi 0.19 nx 1 ny 5 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1 ccov 100
<< end >>
