magic
tech sky130A
magscale 1 2
timestamp 1755691638
<< metal1 >>
rect 25179 2815 25185 3015
rect 25385 2815 26864 3015
rect 26258 2545 26318 2551
rect 26318 2485 26704 2545
rect 26258 2479 26318 2485
rect 26498 1683 26678 2105
rect 29229 1789 29429 2108
rect 26492 1503 26498 1683
rect 26678 1503 26684 1683
rect 29229 1583 29429 1589
rect 25246 1433 25646 1439
rect 25646 1240 25901 1433
rect 25646 1040 26861 1240
rect 25646 1033 25901 1040
rect 25246 1027 25646 1033
<< via1 >>
rect 25185 2815 25385 3015
rect 26258 2485 26318 2545
rect 26498 1503 26678 1683
rect 29229 1589 29429 1789
rect 25246 1033 25646 1433
<< metal2 >>
rect 24099 3015 24299 3024
rect 25185 3015 25385 3021
rect 24299 2815 25185 3015
rect 24099 2806 24299 2815
rect 25185 2809 25385 2815
rect 26143 2545 26199 2552
rect 26141 2543 26258 2545
rect 26141 2487 26143 2543
rect 26199 2487 26258 2543
rect 26141 2485 26258 2487
rect 26318 2485 26324 2545
rect 26143 2478 26199 2485
rect 26498 1683 26678 1689
rect 29223 1589 29229 1789
rect 29429 1589 29435 1789
rect 26498 1443 26678 1503
rect 29229 1493 29429 1589
rect 24821 1433 25211 1437
rect 24816 1428 25246 1433
rect 24816 1038 24821 1428
rect 25211 1038 25246 1428
rect 24816 1033 25246 1038
rect 25646 1033 25652 1433
rect 26494 1273 26503 1443
rect 26673 1273 26682 1443
rect 29229 1284 29429 1293
rect 26498 1268 26678 1273
rect 24821 1029 25211 1033
<< via2 >>
rect 24099 2815 24299 3015
rect 26143 2487 26199 2543
rect 24821 1038 25211 1428
rect 26503 1273 26673 1443
rect 29229 1293 29429 1493
<< metal3 >>
rect 28758 44401 28764 44465
rect 28828 44401 28834 44465
rect 28766 3675 28826 44401
rect 26141 3615 28826 3675
rect 24094 3015 24304 3020
rect 378 2815 384 3015
rect 584 2815 24099 3015
rect 24299 2815 24304 3015
rect 24094 2810 24304 2815
rect 26141 2548 26201 3615
rect 26138 2543 26204 2548
rect 26138 2487 26143 2543
rect 26199 2487 26204 2543
rect 26138 2482 26204 2487
rect 29224 1493 29434 1498
rect 26498 1443 26678 1448
rect 24402 1433 24800 1438
rect 24401 1432 25216 1433
rect 24401 1034 24402 1432
rect 24800 1428 25216 1432
rect 24800 1038 24821 1428
rect 25211 1038 25216 1428
rect 24800 1034 25216 1038
rect 24401 1033 25216 1034
rect 26498 1273 26503 1443
rect 26673 1273 26678 1443
rect 29224 1293 29229 1493
rect 29429 1293 29434 1493
rect 29224 1288 29434 1293
rect 24402 1028 24800 1033
rect 26498 682 26678 1273
rect 29229 1027 29429 1288
rect 29229 821 29429 827
rect 26493 504 26499 682
rect 26677 504 26683 682
rect 26498 503 26678 504
<< via3 >>
rect 28764 44401 28828 44465
rect 384 2815 584 3015
rect 24402 1034 24800 1432
rect 29229 827 29429 1027
rect 26499 504 26677 682
<< metal4 >>
rect 6134 44152 6194 45152
rect 6686 44152 6746 45152
rect 7238 44152 7298 45152
rect 7790 44152 7850 45152
rect 8342 44152 8402 45152
rect 8894 44152 8954 45152
rect 9446 44152 9506 45152
rect 9998 44152 10058 45152
rect 10550 44152 10610 45152
rect 11102 44152 11162 45152
rect 11654 44152 11714 45152
rect 12206 44152 12266 45152
rect 12758 44152 12818 45152
rect 13310 44152 13370 45152
rect 13862 44152 13922 45152
rect 14414 44152 14474 45152
rect 14966 44152 15026 45152
rect 15518 44152 15578 45152
rect 16070 44152 16130 45152
rect 16622 44152 16682 45152
rect 17174 44152 17234 45152
rect 17726 44152 17786 45152
rect 18278 44152 18338 45152
rect 18830 44152 18890 45152
rect 19382 44952 19442 45152
rect 19934 44952 19994 45152
rect 20486 44952 20546 45152
rect 21038 44952 21098 45152
rect 21590 44952 21650 45152
rect 22142 44952 22202 45152
rect 22694 44952 22754 45152
rect 23246 44952 23306 45152
rect 23798 44952 23858 45152
rect 24350 44952 24410 45152
rect 24902 44952 24962 45152
rect 25454 44952 25514 45152
rect 26006 44952 26066 45152
rect 26558 44952 26618 45152
rect 27110 44952 27170 45152
rect 27662 44952 27722 45152
rect 28214 44952 28274 45152
rect 28766 44466 28826 45152
rect 29318 44952 29378 45152
rect 28763 44465 28829 44466
rect 28763 44401 28764 44465
rect 28828 44401 28829 44465
rect 28763 44400 28829 44401
rect 200 3015 600 44152
rect 200 2815 384 3015
rect 584 2815 600 3015
rect 200 1000 600 2815
rect 800 43752 19115 44152
rect 800 1433 1200 43752
rect 800 1432 24801 1433
rect 800 1034 24402 1432
rect 24800 1034 24801 1432
rect 800 1033 24801 1034
rect 800 1000 1200 1033
rect 29228 1027 29430 1028
rect 29228 827 29229 1027
rect 29429 827 29430 1027
rect 29228 826 29430 827
rect 26498 682 26678 683
rect 26498 504 26499 682
rect 26677 504 26678 682
rect 3314 0 3494 200
rect 7178 0 7358 200
rect 11042 0 11222 200
rect 14906 0 15086 200
rect 18770 0 18950 200
rect 22634 0 22814 200
rect 26498 0 26678 504
rect 29229 550 29429 826
rect 30362 550 30542 558
rect 29229 370 30542 550
rect 30362 0 30542 370
use Sample_and_Hold  Sample_and_Hold_0
timestamp 1755657154
transform 1 0 26237 0 1 5645
box 423 -4605 4289 -774
<< labels >>
flabel metal4 s 28766 44952 28826 45152 0 FreeSans 480 90 0 0 clk
port 0 nsew signal input
flabel metal4 s 29318 44952 29378 45152 0 FreeSans 480 90 0 0 ena
port 1 nsew signal input
flabel metal4 s 28214 44952 28274 45152 0 FreeSans 480 90 0 0 rst_n
port 2 nsew signal input
flabel metal4 s 30362 0 30542 200 0 FreeSans 960 0 0 0 ua[0]
port 3 nsew signal bidirectional
flabel metal4 s 26498 0 26678 200 0 FreeSans 960 0 0 0 ua[1]
port 4 nsew signal bidirectional
flabel metal4 s 22634 0 22814 200 0 FreeSans 960 0 0 0 ua[2]
port 5 nsew signal bidirectional
flabel metal4 s 18770 0 18950 200 0 FreeSans 960 0 0 0 ua[3]
port 6 nsew signal bidirectional
flabel metal4 s 14906 0 15086 200 0 FreeSans 960 0 0 0 ua[4]
port 7 nsew signal bidirectional
flabel metal4 s 11042 0 11222 200 0 FreeSans 960 0 0 0 ua[5]
port 8 nsew signal bidirectional
flabel metal4 s 7178 0 7358 200 0 FreeSans 960 0 0 0 ua[6]
port 9 nsew signal bidirectional
flabel metal4 s 3314 0 3494 200 0 FreeSans 960 0 0 0 ua[7]
port 10 nsew signal bidirectional
flabel metal4 s 27662 44952 27722 45152 0 FreeSans 480 90 0 0 ui_in[0]
port 11 nsew signal input
flabel metal4 s 27110 44952 27170 45152 0 FreeSans 480 90 0 0 ui_in[1]
port 12 nsew signal input
flabel metal4 s 26558 44952 26618 45152 0 FreeSans 480 90 0 0 ui_in[2]
port 13 nsew signal input
flabel metal4 s 26006 44952 26066 45152 0 FreeSans 480 90 0 0 ui_in[3]
port 14 nsew signal input
flabel metal4 s 25454 44952 25514 45152 0 FreeSans 480 90 0 0 ui_in[4]
port 15 nsew signal input
flabel metal4 s 24902 44952 24962 45152 0 FreeSans 480 90 0 0 ui_in[5]
port 16 nsew signal input
flabel metal4 s 24350 44952 24410 45152 0 FreeSans 480 90 0 0 ui_in[6]
port 17 nsew signal input
flabel metal4 s 23798 44952 23858 45152 0 FreeSans 480 90 0 0 ui_in[7]
port 18 nsew signal input
flabel metal4 s 23246 44952 23306 45152 0 FreeSans 480 90 0 0 uio_in[0]
port 19 nsew signal input
flabel metal4 s 22694 44952 22754 45152 0 FreeSans 480 90 0 0 uio_in[1]
port 20 nsew signal input
flabel metal4 s 22142 44952 22202 45152 0 FreeSans 480 90 0 0 uio_in[2]
port 21 nsew signal input
flabel metal4 s 21590 44952 21650 45152 0 FreeSans 480 90 0 0 uio_in[3]
port 22 nsew signal input
flabel metal4 s 21038 44952 21098 45152 0 FreeSans 480 90 0 0 uio_in[4]
port 23 nsew signal input
flabel metal4 s 20486 44952 20546 45152 0 FreeSans 480 90 0 0 uio_in[5]
port 24 nsew signal input
flabel metal4 s 19934 44952 19994 45152 0 FreeSans 480 90 0 0 uio_in[6]
port 25 nsew signal input
flabel metal4 s 19382 44952 19442 45152 0 FreeSans 480 90 0 0 uio_in[7]
port 26 nsew signal input
flabel metal4 s 9998 44952 10058 45152 0 FreeSans 480 90 0 0 uio_oe[0]
port 27 nsew signal output
flabel metal4 s 9446 44952 9506 45152 0 FreeSans 480 90 0 0 uio_oe[1]
port 28 nsew signal output
flabel metal4 s 8894 44952 8954 45152 0 FreeSans 480 90 0 0 uio_oe[2]
port 29 nsew signal output
flabel metal4 s 8342 44952 8402 45152 0 FreeSans 480 90 0 0 uio_oe[3]
port 30 nsew signal output
flabel metal4 s 7790 44952 7850 45152 0 FreeSans 480 90 0 0 uio_oe[4]
port 31 nsew signal output
flabel metal4 s 7238 44952 7298 45152 0 FreeSans 480 90 0 0 uio_oe[5]
port 32 nsew signal output
flabel metal4 s 6686 44952 6746 45152 0 FreeSans 480 90 0 0 uio_oe[6]
port 33 nsew signal output
flabel metal4 s 6134 44952 6194 45152 0 FreeSans 480 90 0 0 uio_oe[7]
port 34 nsew signal output
flabel metal4 s 14414 44952 14474 45152 0 FreeSans 480 90 0 0 uio_out[0]
port 35 nsew signal output
flabel metal4 s 13862 44952 13922 45152 0 FreeSans 480 90 0 0 uio_out[1]
port 36 nsew signal output
flabel metal4 s 13310 44952 13370 45152 0 FreeSans 480 90 0 0 uio_out[2]
port 37 nsew signal output
flabel metal4 s 12758 44952 12818 45152 0 FreeSans 480 90 0 0 uio_out[3]
port 38 nsew signal output
flabel metal4 s 12206 44952 12266 45152 0 FreeSans 480 90 0 0 uio_out[4]
port 39 nsew signal output
flabel metal4 s 11654 44952 11714 45152 0 FreeSans 480 90 0 0 uio_out[5]
port 40 nsew signal output
flabel metal4 s 11102 44952 11162 45152 0 FreeSans 480 90 0 0 uio_out[6]
port 41 nsew signal output
flabel metal4 s 10550 44952 10610 45152 0 FreeSans 480 90 0 0 uio_out[7]
port 42 nsew signal output
flabel metal4 s 18830 44952 18890 45152 0 FreeSans 480 90 0 0 uo_out[0]
port 43 nsew signal output
flabel metal4 s 18278 44952 18338 45152 0 FreeSans 480 90 0 0 uo_out[1]
port 44 nsew signal output
flabel metal4 s 17726 44952 17786 45152 0 FreeSans 480 90 0 0 uo_out[2]
port 45 nsew signal output
flabel metal4 s 17174 44952 17234 45152 0 FreeSans 480 90 0 0 uo_out[3]
port 46 nsew signal output
flabel metal4 s 16622 44952 16682 45152 0 FreeSans 480 90 0 0 uo_out[4]
port 47 nsew signal output
flabel metal4 s 16070 44952 16130 45152 0 FreeSans 480 90 0 0 uo_out[5]
port 48 nsew signal output
flabel metal4 s 15518 44952 15578 45152 0 FreeSans 480 90 0 0 uo_out[6]
port 49 nsew signal output
flabel metal4 s 14966 44952 15026 45152 0 FreeSans 480 90 0 0 uo_out[7]
port 50 nsew signal output
flabel metal4 200 1000 600 44152 1 FreeSans 1600 0 0 0 VDPWR
port 51 nsew power bidirectional
flabel metal4 800 1000 1200 44152 1 FreeSans 1600 0 0 0 VGND
port 52 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 32200 45152
<< end >>
