magic
tech sky130A
magscale 1 2
timestamp 1761224974
<< viali >>
rect 2697 15113 2731 15147
rect 8033 14909 8067 14943
rect 8217 14773 8251 14807
rect 15025 14229 15059 14263
rect 9873 13821 9907 13855
rect 9321 13753 9355 13787
rect 9689 13753 9723 13787
rect 10057 13685 10091 13719
rect 10333 13481 10367 13515
rect 11253 13413 11287 13447
rect 8217 13345 8251 13379
rect 10149 13345 10183 13379
rect 8585 13277 8619 13311
rect 10977 13277 11011 13311
rect 12725 13277 12759 13311
rect 13369 13277 13403 13311
rect 10011 13141 10045 13175
rect 12817 13141 12851 13175
rect 15025 13141 15059 13175
rect 8769 12937 8803 12971
rect 10057 12937 10091 12971
rect 9781 12801 9815 12835
rect 10609 12801 10643 12835
rect 11989 12801 12023 12835
rect 8953 12733 8987 12767
rect 9689 12733 9723 12767
rect 10425 12733 10459 12767
rect 11897 12733 11931 12767
rect 15025 12733 15059 12767
rect 9597 12665 9631 12699
rect 10517 12665 10551 12699
rect 9229 12597 9263 12631
rect 12265 12597 12299 12631
rect 13001 12325 13035 12359
rect 7021 12257 7055 12291
rect 10057 12257 10091 12291
rect 7297 12189 7331 12223
rect 10149 12189 10183 12223
rect 12725 12189 12759 12223
rect 14749 12189 14783 12223
rect 10425 12121 10459 12155
rect 8769 12053 8803 12087
rect 7481 11849 7515 11883
rect 12173 11849 12207 11883
rect 10977 11781 11011 11815
rect 11805 11781 11839 11815
rect 15025 11781 15059 11815
rect 9045 11713 9079 11747
rect 10517 11713 10551 11747
rect 7665 11645 7699 11679
rect 8769 11645 8803 11679
rect 10609 11645 10643 11679
rect 11437 11645 11471 11679
rect 11621 11645 11655 11679
rect 11897 11645 11931 11679
rect 12081 11645 12115 11679
rect 12357 11645 12391 11679
rect 12633 11645 12667 11679
rect 12817 11645 12851 11679
rect 12909 11645 12943 11679
rect 13093 11645 13127 11679
rect 11989 11577 12023 11611
rect 8401 11509 8435 11543
rect 8861 11509 8895 11543
rect 13001 11509 13035 11543
rect 10609 11305 10643 11339
rect 11069 11305 11103 11339
rect 11161 11305 11195 11339
rect 12909 11305 12943 11339
rect 9137 11237 9171 11271
rect 13277 11237 13311 11271
rect 6837 11169 6871 11203
rect 9229 11169 9263 11203
rect 9597 11169 9631 11203
rect 10149 11169 10183 11203
rect 10977 11169 11011 11203
rect 12541 11169 12575 11203
rect 7205 11101 7239 11135
rect 8631 11101 8665 11135
rect 9413 11101 9447 11135
rect 10057 11101 10091 11135
rect 11437 11101 11471 11135
rect 12633 11101 12667 11135
rect 13001 11101 13035 11135
rect 15025 11101 15059 11135
rect 8769 10965 8803 10999
rect 9689 10965 9723 10999
rect 10241 10965 10275 10999
rect 7389 10761 7423 10795
rect 10517 10625 10551 10659
rect 15025 10625 15059 10659
rect 7573 10557 7607 10591
rect 10425 10557 10459 10591
rect 10885 10557 10919 10591
rect 11069 10557 11103 10591
rect 12265 10557 12299 10591
rect 12449 10557 12483 10591
rect 10977 10489 11011 10523
rect 10793 10421 10827 10455
rect 12357 10421 12391 10455
rect 12081 10217 12115 10251
rect 12265 10217 12299 10251
rect 11621 10149 11655 10183
rect 11345 10081 11379 10115
rect 11529 10081 11563 10115
rect 11805 10081 11839 10115
rect 11989 10081 12023 10115
rect 12206 10081 12240 10115
rect 12725 10081 12759 10115
rect 13001 10081 13035 10115
rect 6929 10013 6963 10047
rect 7205 10013 7239 10047
rect 12909 10013 12943 10047
rect 11437 9945 11471 9979
rect 8677 9877 8711 9911
rect 12633 9877 12667 9911
rect 13277 9877 13311 9911
rect 15025 9877 15059 9911
rect 7389 9673 7423 9707
rect 12449 9673 12483 9707
rect 12909 9673 12943 9707
rect 8401 9605 8435 9639
rect 8953 9537 8987 9571
rect 7573 9469 7607 9503
rect 9413 9469 9447 9503
rect 9689 9469 9723 9503
rect 12357 9469 12391 9503
rect 12541 9469 12575 9503
rect 12817 9469 12851 9503
rect 13001 9469 13035 9503
rect 15025 9469 15059 9503
rect 11437 9401 11471 9435
rect 8769 9333 8803 9367
rect 8861 9333 8895 9367
rect 9505 9333 9539 9367
rect 8953 9129 8987 9163
rect 12357 9129 12391 9163
rect 10425 9061 10459 9095
rect 13277 9061 13311 9095
rect 6653 8993 6687 9027
rect 7021 8993 7055 9027
rect 9689 8993 9723 9027
rect 9781 8993 9815 9027
rect 10231 8993 10265 9027
rect 10517 8993 10551 9027
rect 12173 8993 12207 9027
rect 12357 8993 12391 9027
rect 13001 8993 13035 9027
rect 8447 8925 8481 8959
rect 9045 8925 9079 8959
rect 9229 8925 9263 8959
rect 10057 8925 10091 8959
rect 10149 8925 10183 8959
rect 15025 8925 15059 8959
rect 10241 8857 10275 8891
rect 8585 8789 8619 8823
rect 9505 8789 9539 8823
rect 7113 8585 7147 8619
rect 11161 8585 11195 8619
rect 9873 8517 9907 8551
rect 10517 8517 10551 8551
rect 11805 8517 11839 8551
rect 9413 8449 9447 8483
rect 10701 8449 10735 8483
rect 10885 8449 10919 8483
rect 11345 8449 11379 8483
rect 12173 8449 12207 8483
rect 7297 8381 7331 8415
rect 9505 8381 9539 8415
rect 10241 8381 10275 8415
rect 10793 8381 10827 8415
rect 10977 8381 11011 8415
rect 11437 8381 11471 8415
rect 12265 8381 12299 8415
rect 15025 8381 15059 8415
rect 10517 8313 10551 8347
rect 10333 8245 10367 8279
rect 12633 8245 12667 8279
rect 8769 8041 8803 8075
rect 10793 8041 10827 8075
rect 11621 8041 11655 8075
rect 15025 7973 15059 8007
rect 7021 7905 7055 7939
rect 9321 7905 9355 7939
rect 11529 7905 11563 7939
rect 11713 7905 11747 7939
rect 12541 7905 12575 7939
rect 13001 7905 13035 7939
rect 7297 7837 7331 7871
rect 9413 7837 9447 7871
rect 9505 7837 9539 7871
rect 10333 7837 10367 7871
rect 10977 7837 11011 7871
rect 11437 7837 11471 7871
rect 12633 7837 12667 7871
rect 12909 7837 12943 7871
rect 13277 7837 13311 7871
rect 10609 7769 10643 7803
rect 11345 7769 11379 7803
rect 8953 7701 8987 7735
rect 7481 7497 7515 7531
rect 12633 7497 12667 7531
rect 13553 7497 13587 7531
rect 14013 7361 14047 7395
rect 7665 7293 7699 7327
rect 9321 7293 9355 7327
rect 11529 7293 11563 7327
rect 12817 7293 12851 7327
rect 13185 7293 13219 7327
rect 13277 7293 13311 7327
rect 13737 7293 13771 7327
rect 13829 7293 13863 7327
rect 13921 7293 13955 7327
rect 9781 7225 9815 7259
rect 12909 7225 12943 7259
rect 13001 7225 13035 7259
rect 9137 7157 9171 7191
rect 10563 6953 10597 6987
rect 12357 6885 12391 6919
rect 9137 6817 9171 6851
rect 11161 6817 11195 6851
rect 11989 6817 12023 6851
rect 12173 6817 12207 6851
rect 12265 6817 12299 6851
rect 12449 6817 12483 6851
rect 12909 6817 12943 6851
rect 6561 6749 6595 6783
rect 6837 6749 6871 6783
rect 8769 6749 8803 6783
rect 11253 6749 11287 6783
rect 11529 6749 11563 6783
rect 8309 6613 8343 6647
rect 12173 6613 12207 6647
rect 13185 6613 13219 6647
rect 13369 6613 13403 6647
rect 7113 6409 7147 6443
rect 8033 6409 8067 6443
rect 9321 6409 9355 6443
rect 8401 6341 8435 6375
rect 9045 6273 9079 6307
rect 9873 6273 9907 6307
rect 13277 6273 13311 6307
rect 13829 6273 13863 6307
rect 7297 6205 7331 6239
rect 9689 6205 9723 6239
rect 9781 6205 9815 6239
rect 13185 6205 13219 6239
rect 13369 6205 13403 6239
rect 13921 6205 13955 6239
rect 8125 6137 8159 6171
rect 8769 6137 8803 6171
rect 8861 6069 8895 6103
rect 13553 6069 13587 6103
rect 9137 5865 9171 5899
rect 8631 5797 8665 5831
rect 9229 5797 9263 5831
rect 13277 5797 13311 5831
rect 6837 5729 6871 5763
rect 9597 5729 9631 5763
rect 7205 5661 7239 5695
rect 9413 5661 9447 5695
rect 10149 5661 10183 5695
rect 13001 5661 13035 5695
rect 15025 5661 15059 5695
rect 9873 5593 9907 5627
rect 10517 5593 10551 5627
rect 8769 5525 8803 5559
rect 10057 5525 10091 5559
rect 10609 5525 10643 5559
rect 7297 5321 7331 5355
rect 11897 5321 11931 5355
rect 13645 5321 13679 5355
rect 11161 5185 11195 5219
rect 12081 5185 12115 5219
rect 12725 5185 12759 5219
rect 7481 5117 7515 5151
rect 9413 5117 9447 5151
rect 11253 5117 11287 5151
rect 11345 5117 11379 5151
rect 11621 5117 11655 5151
rect 11713 5117 11747 5151
rect 12173 5117 12207 5151
rect 12817 5117 12851 5151
rect 13553 5117 13587 5151
rect 13737 5117 13771 5151
rect 11529 5049 11563 5083
rect 12541 4981 12575 5015
rect 13185 4981 13219 5015
rect 10057 4777 10091 4811
rect 10793 4777 10827 4811
rect 10609 4709 10643 4743
rect 12357 4709 12391 4743
rect 9229 4641 9263 4675
rect 9965 4641 9999 4675
rect 10149 4641 10183 4675
rect 10241 4641 10275 4675
rect 11161 4641 11195 4675
rect 11345 4641 11379 4675
rect 11437 4641 11471 4675
rect 12449 4641 12483 4675
rect 13921 4641 13955 4675
rect 11161 4505 11195 4539
rect 9045 4437 9079 4471
rect 10609 4437 10643 4471
rect 13737 4437 13771 4471
rect 8217 4233 8251 4267
rect 13093 4233 13127 4267
rect 13369 4233 13403 4267
rect 14197 4233 14231 4267
rect 10885 4165 10919 4199
rect 11069 4165 11103 4199
rect 11529 4165 11563 4199
rect 13737 4165 13771 4199
rect 6469 4097 6503 4131
rect 8585 4097 8619 4131
rect 8953 4097 8987 4131
rect 10609 4097 10643 4131
rect 11621 4097 11655 4131
rect 11713 4029 11747 4063
rect 11897 4029 11931 4063
rect 13001 4029 13035 4063
rect 13093 4029 13127 4063
rect 13553 4029 13587 4063
rect 13737 4029 13771 4063
rect 13921 4029 13955 4063
rect 14381 4029 14415 4063
rect 14473 4029 14507 4063
rect 6745 3961 6779 3995
rect 11161 3961 11195 3995
rect 10379 3893 10413 3927
rect 11805 3893 11839 3927
rect 7113 3689 7147 3723
rect 8217 3689 8251 3723
rect 9229 3689 9263 3723
rect 9689 3689 9723 3723
rect 12817 3689 12851 3723
rect 8309 3621 8343 3655
rect 9597 3621 9631 3655
rect 13277 3621 13311 3655
rect 7297 3553 7331 3587
rect 8769 3553 8803 3587
rect 9137 3553 9171 3587
rect 11345 3553 11379 3587
rect 12633 3553 12667 3587
rect 13001 3553 13035 3587
rect 8493 3485 8527 3519
rect 9781 3485 9815 3519
rect 11437 3485 11471 3519
rect 11713 3485 11747 3519
rect 12449 3485 12483 3519
rect 15025 3485 15059 3519
rect 7849 3417 7883 3451
rect 6377 3009 6411 3043
rect 12357 3009 12391 3043
rect 9689 2941 9723 2975
rect 12265 2941 12299 2975
rect 6653 2873 6687 2907
rect 8125 2805 8159 2839
rect 9505 2805 9539 2839
rect 12633 2805 12667 2839
rect 7205 2601 7239 2635
rect 8217 2533 8251 2567
rect 7389 2465 7423 2499
rect 8309 2465 8343 2499
rect 8953 2465 8987 2499
rect 9321 2465 9355 2499
rect 12725 2465 12759 2499
rect 13001 2465 13035 2499
rect 15025 2465 15059 2499
rect 8493 2397 8527 2431
rect 12541 2397 12575 2431
rect 13277 2397 13311 2431
rect 7849 2329 7883 2363
rect 10747 2261 10781 2295
rect 12909 2261 12943 2295
rect 9689 2057 9723 2091
rect 11437 2057 11471 2091
rect 13553 2057 13587 2091
rect 11161 1989 11195 2023
rect 8861 1921 8895 1955
rect 9045 1921 9079 1955
rect 10149 1921 10183 1955
rect 10333 1921 10367 1955
rect 11345 1921 11379 1955
rect 12449 1921 12483 1955
rect 8769 1853 8803 1887
rect 11621 1853 11655 1887
rect 11897 1853 11931 1887
rect 11989 1853 12023 1887
rect 12265 1853 12299 1887
rect 12725 1853 12759 1887
rect 13093 1853 13127 1887
rect 13277 1853 13311 1887
rect 13553 1853 13587 1887
rect 13737 1853 13771 1887
rect 10057 1785 10091 1819
rect 10885 1785 10919 1819
rect 8401 1717 8435 1751
rect 11805 1717 11839 1751
rect 12081 1717 12115 1751
rect 12817 1717 12851 1751
rect 13185 1717 13219 1751
rect 8631 1513 8665 1547
rect 12081 1513 12115 1547
rect 15025 1445 15059 1479
rect 6837 1377 6871 1411
rect 8769 1377 8803 1411
rect 11437 1377 11471 1411
rect 13001 1377 13035 1411
rect 7205 1309 7239 1343
rect 9045 1309 9079 1343
rect 11161 1309 11195 1343
rect 12173 1309 12207 1343
rect 13277 1309 13311 1343
rect 10517 1173 10551 1207
rect 12817 1173 12851 1207
rect 7389 969 7423 1003
rect 8585 969 8619 1003
rect 9137 969 9171 1003
rect 11989 969 12023 1003
rect 12449 969 12483 1003
rect 12633 969 12667 1003
rect 12817 969 12851 1003
rect 13185 969 13219 1003
rect 9597 901 9631 935
rect 11897 901 11931 935
rect 10057 833 10091 867
rect 10149 833 10183 867
rect 12081 833 12115 867
rect 12725 833 12759 867
rect 7573 765 7607 799
rect 8401 765 8435 799
rect 9321 765 9355 799
rect 9965 765 9999 799
rect 11805 765 11839 799
rect 12173 765 12207 799
rect 13001 765 13035 799
<< metal1 >>
rect 552 15258 15364 15280
rect 552 15206 2249 15258
rect 2301 15206 2313 15258
rect 2365 15206 2377 15258
rect 2429 15206 2441 15258
rect 2493 15206 2505 15258
rect 2557 15206 5951 15258
rect 6003 15206 6015 15258
rect 6067 15206 6079 15258
rect 6131 15206 6143 15258
rect 6195 15206 6207 15258
rect 6259 15206 9653 15258
rect 9705 15206 9717 15258
rect 9769 15206 9781 15258
rect 9833 15206 9845 15258
rect 9897 15206 9909 15258
rect 9961 15206 13355 15258
rect 13407 15206 13419 15258
rect 13471 15206 13483 15258
rect 13535 15206 13547 15258
rect 13599 15206 13611 15258
rect 13663 15206 15364 15258
rect 552 15184 15364 15206
rect 2682 15104 2688 15156
rect 2740 15104 2746 15156
rect 8018 14900 8024 14952
rect 8076 14900 8082 14952
rect 8202 14764 8208 14816
rect 8260 14764 8266 14816
rect 552 14714 15520 14736
rect 552 14662 4100 14714
rect 4152 14662 4164 14714
rect 4216 14662 4228 14714
rect 4280 14662 4292 14714
rect 4344 14662 4356 14714
rect 4408 14662 7802 14714
rect 7854 14662 7866 14714
rect 7918 14662 7930 14714
rect 7982 14662 7994 14714
rect 8046 14662 8058 14714
rect 8110 14662 11504 14714
rect 11556 14662 11568 14714
rect 11620 14662 11632 14714
rect 11684 14662 11696 14714
rect 11748 14662 11760 14714
rect 11812 14662 15206 14714
rect 15258 14662 15270 14714
rect 15322 14662 15334 14714
rect 15386 14662 15398 14714
rect 15450 14662 15462 14714
rect 15514 14662 15520 14714
rect 552 14640 15520 14662
rect 15010 14220 15016 14272
rect 15068 14220 15074 14272
rect 552 14170 15364 14192
rect 552 14118 2249 14170
rect 2301 14118 2313 14170
rect 2365 14118 2377 14170
rect 2429 14118 2441 14170
rect 2493 14118 2505 14170
rect 2557 14118 5951 14170
rect 6003 14118 6015 14170
rect 6067 14118 6079 14170
rect 6131 14118 6143 14170
rect 6195 14118 6207 14170
rect 6259 14118 9653 14170
rect 9705 14118 9717 14170
rect 9769 14118 9781 14170
rect 9833 14118 9845 14170
rect 9897 14118 9909 14170
rect 9961 14118 13355 14170
rect 13407 14118 13419 14170
rect 13471 14118 13483 14170
rect 13535 14118 13547 14170
rect 13599 14118 13611 14170
rect 13663 14118 15364 14170
rect 552 14096 15364 14118
rect 8202 13812 8208 13864
rect 8260 13852 8266 13864
rect 9861 13855 9919 13861
rect 9861 13852 9873 13855
rect 8260 13824 9873 13852
rect 8260 13812 8266 13824
rect 9861 13821 9873 13824
rect 9907 13821 9919 13855
rect 9861 13815 9919 13821
rect 8662 13744 8668 13796
rect 8720 13784 8726 13796
rect 9309 13787 9367 13793
rect 9309 13784 9321 13787
rect 8720 13756 9321 13784
rect 8720 13744 8726 13756
rect 9309 13753 9321 13756
rect 9355 13753 9367 13787
rect 9309 13747 9367 13753
rect 9677 13787 9735 13793
rect 9677 13753 9689 13787
rect 9723 13784 9735 13787
rect 9723 13756 10088 13784
rect 9723 13753 9735 13756
rect 9677 13747 9735 13753
rect 10060 13725 10088 13756
rect 10045 13719 10103 13725
rect 10045 13685 10057 13719
rect 10091 13716 10103 13719
rect 11882 13716 11888 13728
rect 10091 13688 11888 13716
rect 10091 13685 10103 13688
rect 10045 13679 10103 13685
rect 11882 13676 11888 13688
rect 11940 13676 11946 13728
rect 552 13626 15520 13648
rect 552 13574 4100 13626
rect 4152 13574 4164 13626
rect 4216 13574 4228 13626
rect 4280 13574 4292 13626
rect 4344 13574 4356 13626
rect 4408 13574 7802 13626
rect 7854 13574 7866 13626
rect 7918 13574 7930 13626
rect 7982 13574 7994 13626
rect 8046 13574 8058 13626
rect 8110 13574 11504 13626
rect 11556 13574 11568 13626
rect 11620 13574 11632 13626
rect 11684 13574 11696 13626
rect 11748 13574 11760 13626
rect 11812 13574 15206 13626
rect 15258 13574 15270 13626
rect 15322 13574 15334 13626
rect 15386 13574 15398 13626
rect 15450 13574 15462 13626
rect 15514 13574 15520 13626
rect 552 13552 15520 13574
rect 8662 13472 8668 13524
rect 8720 13512 8726 13524
rect 10321 13515 10379 13521
rect 8720 13484 8892 13512
rect 8720 13472 8726 13484
rect 8864 13444 8892 13484
rect 10321 13481 10333 13515
rect 10367 13512 10379 13515
rect 10367 13484 11284 13512
rect 10367 13481 10379 13484
rect 10321 13475 10379 13481
rect 11256 13453 11284 13484
rect 11241 13447 11299 13453
rect 8864 13416 8970 13444
rect 11241 13413 11253 13447
rect 11287 13413 11299 13447
rect 11241 13407 11299 13413
rect 11882 13404 11888 13456
rect 11940 13404 11946 13456
rect 7006 13336 7012 13388
rect 7064 13376 7070 13388
rect 8205 13379 8263 13385
rect 8205 13376 8217 13379
rect 7064 13348 8217 13376
rect 7064 13336 7070 13348
rect 8205 13345 8217 13348
rect 8251 13376 8263 13379
rect 8251 13348 8708 13376
rect 8251 13345 8263 13348
rect 8205 13339 8263 13345
rect 8570 13268 8576 13320
rect 8628 13268 8634 13320
rect 8680 13308 8708 13348
rect 10134 13336 10140 13388
rect 10192 13336 10198 13388
rect 10962 13308 10968 13320
rect 8680 13280 10968 13308
rect 10962 13268 10968 13280
rect 11020 13268 11026 13320
rect 11238 13268 11244 13320
rect 11296 13308 11302 13320
rect 12713 13311 12771 13317
rect 12713 13308 12725 13311
rect 11296 13280 12725 13308
rect 11296 13268 11302 13280
rect 12713 13277 12725 13280
rect 12759 13308 12771 13311
rect 13357 13311 13415 13317
rect 13357 13308 13369 13311
rect 12759 13280 13369 13308
rect 12759 13277 12771 13280
rect 12713 13271 12771 13277
rect 13357 13277 13369 13280
rect 13403 13277 13415 13311
rect 13357 13271 13415 13277
rect 10042 13181 10048 13184
rect 9999 13175 10048 13181
rect 9999 13141 10011 13175
rect 10045 13141 10048 13175
rect 9999 13135 10048 13141
rect 10042 13132 10048 13135
rect 10100 13132 10106 13184
rect 12802 13132 12808 13184
rect 12860 13132 12866 13184
rect 15010 13132 15016 13184
rect 15068 13132 15074 13184
rect 552 13082 15364 13104
rect 552 13030 2249 13082
rect 2301 13030 2313 13082
rect 2365 13030 2377 13082
rect 2429 13030 2441 13082
rect 2493 13030 2505 13082
rect 2557 13030 5951 13082
rect 6003 13030 6015 13082
rect 6067 13030 6079 13082
rect 6131 13030 6143 13082
rect 6195 13030 6207 13082
rect 6259 13030 9653 13082
rect 9705 13030 9717 13082
rect 9769 13030 9781 13082
rect 9833 13030 9845 13082
rect 9897 13030 9909 13082
rect 9961 13030 13355 13082
rect 13407 13030 13419 13082
rect 13471 13030 13483 13082
rect 13535 13030 13547 13082
rect 13599 13030 13611 13082
rect 13663 13030 15364 13082
rect 552 13008 15364 13030
rect 8570 12928 8576 12980
rect 8628 12968 8634 12980
rect 8757 12971 8815 12977
rect 8757 12968 8769 12971
rect 8628 12940 8769 12968
rect 8628 12928 8634 12940
rect 8757 12937 8769 12940
rect 8803 12937 8815 12971
rect 8757 12931 8815 12937
rect 10045 12971 10103 12977
rect 10045 12937 10057 12971
rect 10091 12968 10103 12971
rect 10134 12968 10140 12980
rect 10091 12940 10140 12968
rect 10091 12937 10103 12940
rect 10045 12931 10103 12937
rect 10134 12928 10140 12940
rect 10192 12928 10198 12980
rect 9398 12792 9404 12844
rect 9456 12832 9462 12844
rect 9769 12835 9827 12841
rect 9769 12832 9781 12835
rect 9456 12804 9781 12832
rect 9456 12792 9462 12804
rect 9769 12801 9781 12804
rect 9815 12801 9827 12835
rect 9769 12795 9827 12801
rect 10226 12792 10232 12844
rect 10284 12832 10290 12844
rect 10597 12835 10655 12841
rect 10597 12832 10609 12835
rect 10284 12804 10609 12832
rect 10284 12792 10290 12804
rect 10597 12801 10609 12804
rect 10643 12801 10655 12835
rect 10597 12795 10655 12801
rect 11974 12792 11980 12844
rect 12032 12792 12038 12844
rect 8941 12767 8999 12773
rect 8941 12733 8953 12767
rect 8987 12764 8999 12767
rect 9677 12767 9735 12773
rect 8987 12736 9260 12764
rect 8987 12733 8999 12736
rect 8941 12727 8999 12733
rect 9232 12637 9260 12736
rect 9677 12733 9689 12767
rect 9723 12764 9735 12767
rect 10042 12764 10048 12776
rect 9723 12736 10048 12764
rect 9723 12733 9735 12736
rect 9677 12727 9735 12733
rect 10042 12724 10048 12736
rect 10100 12724 10106 12776
rect 10134 12724 10140 12776
rect 10192 12764 10198 12776
rect 10413 12767 10471 12773
rect 10413 12764 10425 12767
rect 10192 12736 10425 12764
rect 10192 12724 10198 12736
rect 10413 12733 10425 12736
rect 10459 12764 10471 12767
rect 11238 12764 11244 12776
rect 10459 12736 11244 12764
rect 10459 12733 10471 12736
rect 10413 12727 10471 12733
rect 11238 12724 11244 12736
rect 11296 12724 11302 12776
rect 11885 12767 11943 12773
rect 11885 12733 11897 12767
rect 11931 12764 11943 12767
rect 12802 12764 12808 12776
rect 11931 12736 12808 12764
rect 11931 12733 11943 12736
rect 11885 12727 11943 12733
rect 12802 12724 12808 12736
rect 12860 12724 12866 12776
rect 15010 12724 15016 12776
rect 15068 12724 15074 12776
rect 9585 12699 9643 12705
rect 9585 12665 9597 12699
rect 9631 12696 9643 12699
rect 10505 12699 10563 12705
rect 10505 12696 10517 12699
rect 9631 12668 10517 12696
rect 9631 12665 9643 12668
rect 9585 12659 9643 12665
rect 10505 12665 10517 12668
rect 10551 12696 10563 12699
rect 14734 12696 14740 12708
rect 10551 12668 14740 12696
rect 10551 12665 10563 12668
rect 10505 12659 10563 12665
rect 14734 12656 14740 12668
rect 14792 12656 14798 12708
rect 9217 12631 9275 12637
rect 9217 12597 9229 12631
rect 9263 12597 9275 12631
rect 9217 12591 9275 12597
rect 12250 12588 12256 12640
rect 12308 12588 12314 12640
rect 552 12538 15520 12560
rect 552 12486 4100 12538
rect 4152 12486 4164 12538
rect 4216 12486 4228 12538
rect 4280 12486 4292 12538
rect 4344 12486 4356 12538
rect 4408 12486 7802 12538
rect 7854 12486 7866 12538
rect 7918 12486 7930 12538
rect 7982 12486 7994 12538
rect 8046 12486 8058 12538
rect 8110 12486 11504 12538
rect 11556 12486 11568 12538
rect 11620 12486 11632 12538
rect 11684 12486 11696 12538
rect 11748 12486 11760 12538
rect 11812 12486 15206 12538
rect 15258 12486 15270 12538
rect 15322 12486 15334 12538
rect 15386 12486 15398 12538
rect 15450 12486 15462 12538
rect 15514 12486 15520 12538
rect 552 12464 15520 12486
rect 8662 12356 8668 12368
rect 8510 12328 8668 12356
rect 8662 12316 8668 12328
rect 8720 12316 8726 12368
rect 12250 12316 12256 12368
rect 12308 12356 12314 12368
rect 12989 12359 13047 12365
rect 12989 12356 13001 12359
rect 12308 12328 13001 12356
rect 12308 12316 12314 12328
rect 12989 12325 13001 12328
rect 13035 12325 13047 12359
rect 12989 12319 13047 12325
rect 7006 12248 7012 12300
rect 7064 12248 7070 12300
rect 10042 12248 10048 12300
rect 10100 12248 10106 12300
rect 7282 12180 7288 12232
rect 7340 12180 7346 12232
rect 10134 12180 10140 12232
rect 10192 12180 10198 12232
rect 10962 12180 10968 12232
rect 11020 12220 11026 12232
rect 12713 12223 12771 12229
rect 12713 12220 12725 12223
rect 11020 12192 12725 12220
rect 11020 12180 11026 12192
rect 12713 12189 12725 12192
rect 12759 12189 12771 12223
rect 12713 12183 12771 12189
rect 10413 12155 10471 12161
rect 10413 12121 10425 12155
rect 10459 12152 10471 12155
rect 10502 12152 10508 12164
rect 10459 12124 10508 12152
rect 10459 12121 10471 12124
rect 10413 12115 10471 12121
rect 10502 12112 10508 12124
rect 10560 12112 10566 12164
rect 8754 12044 8760 12096
rect 8812 12044 8818 12096
rect 12728 12084 12756 12183
rect 13722 12180 13728 12232
rect 13780 12220 13786 12232
rect 14108 12220 14136 12274
rect 13780 12192 14136 12220
rect 13780 12180 13786 12192
rect 14734 12180 14740 12232
rect 14792 12180 14798 12232
rect 12986 12084 12992 12096
rect 12728 12056 12992 12084
rect 12986 12044 12992 12056
rect 13044 12044 13050 12096
rect 552 11994 15364 12016
rect 552 11942 2249 11994
rect 2301 11942 2313 11994
rect 2365 11942 2377 11994
rect 2429 11942 2441 11994
rect 2493 11942 2505 11994
rect 2557 11942 5951 11994
rect 6003 11942 6015 11994
rect 6067 11942 6079 11994
rect 6131 11942 6143 11994
rect 6195 11942 6207 11994
rect 6259 11942 9653 11994
rect 9705 11942 9717 11994
rect 9769 11942 9781 11994
rect 9833 11942 9845 11994
rect 9897 11942 9909 11994
rect 9961 11942 13355 11994
rect 13407 11942 13419 11994
rect 13471 11942 13483 11994
rect 13535 11942 13547 11994
rect 13599 11942 13611 11994
rect 13663 11942 15364 11994
rect 552 11920 15364 11942
rect 7282 11840 7288 11892
rect 7340 11880 7346 11892
rect 7469 11883 7527 11889
rect 7469 11880 7481 11883
rect 7340 11852 7481 11880
rect 7340 11840 7346 11852
rect 7469 11849 7481 11852
rect 7515 11849 7527 11883
rect 7469 11843 7527 11849
rect 11974 11840 11980 11892
rect 12032 11880 12038 11892
rect 12161 11883 12219 11889
rect 12161 11880 12173 11883
rect 12032 11852 12173 11880
rect 12032 11840 12038 11852
rect 12161 11849 12173 11852
rect 12207 11849 12219 11883
rect 12161 11843 12219 11849
rect 10965 11815 11023 11821
rect 10965 11781 10977 11815
rect 11011 11781 11023 11815
rect 10965 11775 11023 11781
rect 11793 11815 11851 11821
rect 11793 11781 11805 11815
rect 11839 11812 11851 11815
rect 15013 11815 15071 11821
rect 11839 11784 12388 11812
rect 11839 11781 11851 11784
rect 11793 11775 11851 11781
rect 8938 11704 8944 11756
rect 8996 11744 9002 11756
rect 9033 11747 9091 11753
rect 9033 11744 9045 11747
rect 8996 11716 9045 11744
rect 8996 11704 9002 11716
rect 9033 11713 9045 11716
rect 9079 11744 9091 11747
rect 10226 11744 10232 11756
rect 9079 11716 10232 11744
rect 9079 11713 9091 11716
rect 9033 11707 9091 11713
rect 10226 11704 10232 11716
rect 10284 11704 10290 11756
rect 10502 11704 10508 11756
rect 10560 11704 10566 11756
rect 10980 11744 11008 11775
rect 12360 11744 12388 11784
rect 15013 11781 15025 11815
rect 15059 11812 15071 11815
rect 15654 11812 15660 11824
rect 15059 11784 15660 11812
rect 15059 11781 15071 11784
rect 15013 11775 15071 11781
rect 15654 11772 15660 11784
rect 15712 11772 15718 11824
rect 10980 11716 12112 11744
rect 7653 11679 7711 11685
rect 7653 11645 7665 11679
rect 7699 11676 7711 11679
rect 7699 11648 8432 11676
rect 7699 11645 7711 11648
rect 7653 11639 7711 11645
rect 8404 11549 8432 11648
rect 8754 11636 8760 11688
rect 8812 11636 8818 11688
rect 10597 11679 10655 11685
rect 10597 11645 10609 11679
rect 10643 11676 10655 11679
rect 11146 11676 11152 11688
rect 10643 11648 11152 11676
rect 10643 11645 10655 11648
rect 10597 11639 10655 11645
rect 11146 11636 11152 11648
rect 11204 11636 11210 11688
rect 11624 11685 11652 11716
rect 12084 11685 12112 11716
rect 12360 11716 13124 11744
rect 12360 11685 12388 11716
rect 11425 11679 11483 11685
rect 11425 11645 11437 11679
rect 11471 11645 11483 11679
rect 11425 11639 11483 11645
rect 11609 11679 11667 11685
rect 11609 11645 11621 11679
rect 11655 11645 11667 11679
rect 11609 11639 11667 11645
rect 11885 11679 11943 11685
rect 11885 11645 11897 11679
rect 11931 11645 11943 11679
rect 11885 11639 11943 11645
rect 12069 11679 12127 11685
rect 12069 11645 12081 11679
rect 12115 11645 12127 11679
rect 12069 11639 12127 11645
rect 12345 11679 12403 11685
rect 12345 11645 12357 11679
rect 12391 11645 12403 11679
rect 12345 11639 12403 11645
rect 12621 11679 12679 11685
rect 12621 11645 12633 11679
rect 12667 11645 12679 11679
rect 12621 11639 12679 11645
rect 10134 11568 10140 11620
rect 10192 11608 10198 11620
rect 11440 11608 11468 11639
rect 11900 11608 11928 11639
rect 10192 11580 11928 11608
rect 11977 11611 12035 11617
rect 10192 11568 10198 11580
rect 11977 11577 11989 11611
rect 12023 11608 12035 11611
rect 12636 11608 12664 11639
rect 12802 11636 12808 11688
rect 12860 11636 12866 11688
rect 13096 11685 13124 11716
rect 12897 11679 12955 11685
rect 12897 11645 12909 11679
rect 12943 11645 12955 11679
rect 12897 11639 12955 11645
rect 13081 11679 13139 11685
rect 13081 11645 13093 11679
rect 13127 11645 13139 11679
rect 13081 11639 13139 11645
rect 12912 11608 12940 11639
rect 12023 11580 12940 11608
rect 12023 11577 12035 11580
rect 11977 11571 12035 11577
rect 8389 11543 8447 11549
rect 8389 11509 8401 11543
rect 8435 11509 8447 11543
rect 8389 11503 8447 11509
rect 8846 11500 8852 11552
rect 8904 11500 8910 11552
rect 12618 11500 12624 11552
rect 12676 11540 12682 11552
rect 12989 11543 13047 11549
rect 12989 11540 13001 11543
rect 12676 11512 13001 11540
rect 12676 11500 12682 11512
rect 12989 11509 13001 11512
rect 13035 11509 13047 11543
rect 12989 11503 13047 11509
rect 552 11450 15520 11472
rect 552 11398 4100 11450
rect 4152 11398 4164 11450
rect 4216 11398 4228 11450
rect 4280 11398 4292 11450
rect 4344 11398 4356 11450
rect 4408 11398 7802 11450
rect 7854 11398 7866 11450
rect 7918 11398 7930 11450
rect 7982 11398 7994 11450
rect 8046 11398 8058 11450
rect 8110 11398 11504 11450
rect 11556 11398 11568 11450
rect 11620 11398 11632 11450
rect 11684 11398 11696 11450
rect 11748 11398 11760 11450
rect 11812 11398 15206 11450
rect 15258 11398 15270 11450
rect 15322 11398 15334 11450
rect 15386 11398 15398 11450
rect 15450 11398 15462 11450
rect 15514 11398 15520 11450
rect 552 11376 15520 11398
rect 10597 11339 10655 11345
rect 10597 11305 10609 11339
rect 10643 11336 10655 11339
rect 10870 11336 10876 11348
rect 10643 11308 10876 11336
rect 10643 11305 10655 11308
rect 10597 11299 10655 11305
rect 10870 11296 10876 11308
rect 10928 11336 10934 11348
rect 11057 11339 11115 11345
rect 11057 11336 11069 11339
rect 10928 11308 11069 11336
rect 10928 11296 10934 11308
rect 11057 11305 11069 11308
rect 11103 11305 11115 11339
rect 11057 11299 11115 11305
rect 11146 11296 11152 11348
rect 11204 11296 11210 11348
rect 12897 11339 12955 11345
rect 12897 11305 12909 11339
rect 12943 11305 12955 11339
rect 12897 11299 12955 11305
rect 8662 11268 8668 11280
rect 8234 11240 8668 11268
rect 8662 11228 8668 11240
rect 8720 11228 8726 11280
rect 8846 11228 8852 11280
rect 8904 11268 8910 11280
rect 9125 11271 9183 11277
rect 9125 11268 9137 11271
rect 8904 11240 9137 11268
rect 8904 11228 8910 11240
rect 9125 11237 9137 11240
rect 9171 11268 9183 11271
rect 12912 11268 12940 11299
rect 13265 11271 13323 11277
rect 13265 11268 13277 11271
rect 9171 11240 12020 11268
rect 12912 11240 13277 11268
rect 9171 11237 9183 11240
rect 9125 11231 9183 11237
rect 6825 11203 6883 11209
rect 6825 11169 6837 11203
rect 6871 11200 6883 11203
rect 6914 11200 6920 11212
rect 6871 11172 6920 11200
rect 6871 11169 6883 11172
rect 6825 11163 6883 11169
rect 6914 11160 6920 11172
rect 6972 11160 6978 11212
rect 9217 11203 9275 11209
rect 9217 11169 9229 11203
rect 9263 11200 9275 11203
rect 9585 11203 9643 11209
rect 9585 11200 9597 11203
rect 9263 11172 9597 11200
rect 9263 11169 9275 11172
rect 9217 11163 9275 11169
rect 9585 11169 9597 11172
rect 9631 11169 9643 11203
rect 9585 11163 9643 11169
rect 7190 11092 7196 11144
rect 7248 11092 7254 11144
rect 8619 11135 8677 11141
rect 8619 11101 8631 11135
rect 8665 11132 8677 11135
rect 9232 11132 9260 11163
rect 8665 11104 9260 11132
rect 8665 11101 8677 11104
rect 8619 11095 8677 11101
rect 9398 11092 9404 11144
rect 9456 11092 9462 11144
rect 9600 11064 9628 11163
rect 10134 11160 10140 11212
rect 10192 11160 10198 11212
rect 10965 11203 11023 11209
rect 10965 11169 10977 11203
rect 11011 11200 11023 11203
rect 11146 11200 11152 11212
rect 11011 11172 11152 11200
rect 11011 11169 11023 11172
rect 10965 11163 11023 11169
rect 11146 11160 11152 11172
rect 11204 11160 11210 11212
rect 10045 11135 10103 11141
rect 10045 11101 10057 11135
rect 10091 11132 10103 11135
rect 11054 11132 11060 11144
rect 10091 11104 11060 11132
rect 10091 11101 10103 11104
rect 10045 11095 10103 11101
rect 11054 11092 11060 11104
rect 11112 11132 11118 11144
rect 11425 11135 11483 11141
rect 11425 11132 11437 11135
rect 11112 11104 11437 11132
rect 11112 11092 11118 11104
rect 11425 11101 11437 11104
rect 11471 11101 11483 11135
rect 11425 11095 11483 11101
rect 11992 11064 12020 11240
rect 13265 11237 13277 11240
rect 13311 11237 13323 11271
rect 13265 11231 13323 11237
rect 13722 11228 13728 11280
rect 13780 11228 13786 11280
rect 12066 11160 12072 11212
rect 12124 11200 12130 11212
rect 12529 11203 12587 11209
rect 12529 11200 12541 11203
rect 12124 11172 12541 11200
rect 12124 11160 12130 11172
rect 12529 11169 12541 11172
rect 12575 11200 12587 11203
rect 12802 11200 12808 11212
rect 12575 11172 12808 11200
rect 12575 11169 12587 11172
rect 12529 11163 12587 11169
rect 12802 11160 12808 11172
rect 12860 11160 12866 11212
rect 12618 11092 12624 11144
rect 12676 11092 12682 11144
rect 12986 11092 12992 11144
rect 13044 11092 13050 11144
rect 14918 11132 14924 11144
rect 13096 11104 14924 11132
rect 13096 11064 13124 11104
rect 14918 11092 14924 11104
rect 14976 11132 14982 11144
rect 15013 11135 15071 11141
rect 15013 11132 15025 11135
rect 14976 11104 15025 11132
rect 14976 11092 14982 11104
rect 15013 11101 15025 11104
rect 15059 11101 15071 11135
rect 15013 11095 15071 11101
rect 9600 11036 10272 11064
rect 11992 11036 13124 11064
rect 8754 10956 8760 11008
rect 8812 10956 8818 11008
rect 8846 10956 8852 11008
rect 8904 10996 8910 11008
rect 9677 10999 9735 11005
rect 9677 10996 9689 10999
rect 8904 10968 9689 10996
rect 8904 10956 8910 10968
rect 9677 10965 9689 10968
rect 9723 10996 9735 10999
rect 10134 10996 10140 11008
rect 9723 10968 10140 10996
rect 9723 10965 9735 10968
rect 9677 10959 9735 10965
rect 10134 10956 10140 10968
rect 10192 10956 10198 11008
rect 10244 11005 10272 11036
rect 10229 10999 10287 11005
rect 10229 10965 10241 10999
rect 10275 10965 10287 10999
rect 10229 10959 10287 10965
rect 552 10906 15364 10928
rect 552 10854 2249 10906
rect 2301 10854 2313 10906
rect 2365 10854 2377 10906
rect 2429 10854 2441 10906
rect 2493 10854 2505 10906
rect 2557 10854 5951 10906
rect 6003 10854 6015 10906
rect 6067 10854 6079 10906
rect 6131 10854 6143 10906
rect 6195 10854 6207 10906
rect 6259 10854 9653 10906
rect 9705 10854 9717 10906
rect 9769 10854 9781 10906
rect 9833 10854 9845 10906
rect 9897 10854 9909 10906
rect 9961 10854 13355 10906
rect 13407 10854 13419 10906
rect 13471 10854 13483 10906
rect 13535 10854 13547 10906
rect 13599 10854 13611 10906
rect 13663 10854 15364 10906
rect 552 10832 15364 10854
rect 7190 10752 7196 10804
rect 7248 10792 7254 10804
rect 7377 10795 7435 10801
rect 7377 10792 7389 10795
rect 7248 10764 7389 10792
rect 7248 10752 7254 10764
rect 7377 10761 7389 10764
rect 7423 10761 7435 10795
rect 7377 10755 7435 10761
rect 10505 10659 10563 10665
rect 10505 10625 10517 10659
rect 10551 10656 10563 10659
rect 11146 10656 11152 10668
rect 10551 10628 11152 10656
rect 10551 10625 10563 10628
rect 10505 10619 10563 10625
rect 11146 10616 11152 10628
rect 11204 10616 11210 10668
rect 15010 10616 15016 10668
rect 15068 10616 15074 10668
rect 7561 10591 7619 10597
rect 7561 10557 7573 10591
rect 7607 10588 7619 10591
rect 8754 10588 8760 10600
rect 7607 10560 8760 10588
rect 7607 10557 7619 10560
rect 7561 10551 7619 10557
rect 8754 10548 8760 10560
rect 8812 10548 8818 10600
rect 10413 10591 10471 10597
rect 10413 10557 10425 10591
rect 10459 10557 10471 10591
rect 10413 10551 10471 10557
rect 10428 10520 10456 10551
rect 10870 10548 10876 10600
rect 10928 10548 10934 10600
rect 11054 10548 11060 10600
rect 11112 10548 11118 10600
rect 11974 10548 11980 10600
rect 12032 10588 12038 10600
rect 12253 10591 12311 10597
rect 12253 10588 12265 10591
rect 12032 10560 12265 10588
rect 12032 10548 12038 10560
rect 12253 10557 12265 10560
rect 12299 10557 12311 10591
rect 12253 10551 12311 10557
rect 12434 10548 12440 10600
rect 12492 10548 12498 10600
rect 10965 10523 11023 10529
rect 10965 10520 10977 10523
rect 10428 10492 10977 10520
rect 10965 10489 10977 10492
rect 11011 10489 11023 10523
rect 10965 10483 11023 10489
rect 10781 10455 10839 10461
rect 10781 10421 10793 10455
rect 10827 10452 10839 10455
rect 11330 10452 11336 10464
rect 10827 10424 11336 10452
rect 10827 10421 10839 10424
rect 10781 10415 10839 10421
rect 11330 10412 11336 10424
rect 11388 10412 11394 10464
rect 12342 10412 12348 10464
rect 12400 10412 12406 10464
rect 552 10362 15520 10384
rect 552 10310 4100 10362
rect 4152 10310 4164 10362
rect 4216 10310 4228 10362
rect 4280 10310 4292 10362
rect 4344 10310 4356 10362
rect 4408 10310 7802 10362
rect 7854 10310 7866 10362
rect 7918 10310 7930 10362
rect 7982 10310 7994 10362
rect 8046 10310 8058 10362
rect 8110 10310 11504 10362
rect 11556 10310 11568 10362
rect 11620 10310 11632 10362
rect 11684 10310 11696 10362
rect 11748 10310 11760 10362
rect 11812 10310 15206 10362
rect 15258 10310 15270 10362
rect 15322 10310 15334 10362
rect 15386 10310 15398 10362
rect 15450 10310 15462 10362
rect 15514 10310 15520 10362
rect 552 10288 15520 10310
rect 12066 10208 12072 10260
rect 12124 10208 12130 10260
rect 12250 10208 12256 10260
rect 12308 10208 12314 10260
rect 8662 10180 8668 10192
rect 8418 10152 8668 10180
rect 8662 10140 8668 10152
rect 8720 10140 8726 10192
rect 11609 10183 11667 10189
rect 11609 10180 11621 10183
rect 11348 10152 11621 10180
rect 11348 10124 11376 10152
rect 11609 10149 11621 10152
rect 11655 10149 11667 10183
rect 11609 10143 11667 10149
rect 11330 10072 11336 10124
rect 11388 10072 11394 10124
rect 11422 10072 11428 10124
rect 11480 10112 11486 10124
rect 11517 10115 11575 10121
rect 11517 10112 11529 10115
rect 11480 10084 11529 10112
rect 11480 10072 11486 10084
rect 11517 10081 11529 10084
rect 11563 10112 11575 10115
rect 11793 10115 11851 10121
rect 11793 10112 11805 10115
rect 11563 10084 11805 10112
rect 11563 10081 11575 10084
rect 11517 10075 11575 10081
rect 11793 10081 11805 10084
rect 11839 10081 11851 10115
rect 11793 10075 11851 10081
rect 11974 10072 11980 10124
rect 12032 10112 12038 10124
rect 12194 10115 12252 10121
rect 12194 10112 12206 10115
rect 12032 10084 12206 10112
rect 12032 10072 12038 10084
rect 12194 10081 12206 10084
rect 12240 10081 12252 10115
rect 12194 10075 12252 10081
rect 12342 10072 12348 10124
rect 12400 10112 12406 10124
rect 12713 10115 12771 10121
rect 12713 10112 12725 10115
rect 12400 10084 12725 10112
rect 12400 10072 12406 10084
rect 12713 10081 12725 10084
rect 12759 10112 12771 10115
rect 12989 10115 13047 10121
rect 12989 10112 13001 10115
rect 12759 10084 13001 10112
rect 12759 10081 12771 10084
rect 12713 10075 12771 10081
rect 12989 10081 13001 10084
rect 13035 10081 13047 10115
rect 12989 10075 13047 10081
rect 6914 10004 6920 10056
rect 6972 10004 6978 10056
rect 7190 10004 7196 10056
rect 7248 10004 7254 10056
rect 12894 10004 12900 10056
rect 12952 10004 12958 10056
rect 11425 9979 11483 9985
rect 11425 9945 11437 9979
rect 11471 9976 11483 9979
rect 12434 9976 12440 9988
rect 11471 9948 12440 9976
rect 11471 9945 11483 9948
rect 11425 9939 11483 9945
rect 12434 9936 12440 9948
rect 12492 9936 12498 9988
rect 8665 9911 8723 9917
rect 8665 9877 8677 9911
rect 8711 9908 8723 9911
rect 8754 9908 8760 9920
rect 8711 9880 8760 9908
rect 8711 9877 8723 9880
rect 8665 9871 8723 9877
rect 8754 9868 8760 9880
rect 8812 9868 8818 9920
rect 12621 9911 12679 9917
rect 12621 9877 12633 9911
rect 12667 9908 12679 9911
rect 12802 9908 12808 9920
rect 12667 9880 12808 9908
rect 12667 9877 12679 9880
rect 12621 9871 12679 9877
rect 12802 9868 12808 9880
rect 12860 9868 12866 9920
rect 13170 9868 13176 9920
rect 13228 9908 13234 9920
rect 13265 9911 13323 9917
rect 13265 9908 13277 9911
rect 13228 9880 13277 9908
rect 13228 9868 13234 9880
rect 13265 9877 13277 9880
rect 13311 9877 13323 9911
rect 13265 9871 13323 9877
rect 15010 9868 15016 9920
rect 15068 9868 15074 9920
rect 552 9818 15364 9840
rect 552 9766 2249 9818
rect 2301 9766 2313 9818
rect 2365 9766 2377 9818
rect 2429 9766 2441 9818
rect 2493 9766 2505 9818
rect 2557 9766 5951 9818
rect 6003 9766 6015 9818
rect 6067 9766 6079 9818
rect 6131 9766 6143 9818
rect 6195 9766 6207 9818
rect 6259 9766 9653 9818
rect 9705 9766 9717 9818
rect 9769 9766 9781 9818
rect 9833 9766 9845 9818
rect 9897 9766 9909 9818
rect 9961 9766 13355 9818
rect 13407 9766 13419 9818
rect 13471 9766 13483 9818
rect 13535 9766 13547 9818
rect 13599 9766 13611 9818
rect 13663 9766 15364 9818
rect 552 9744 15364 9766
rect 7190 9664 7196 9716
rect 7248 9704 7254 9716
rect 7377 9707 7435 9713
rect 7377 9704 7389 9707
rect 7248 9676 7389 9704
rect 7248 9664 7254 9676
rect 7377 9673 7389 9676
rect 7423 9673 7435 9707
rect 7377 9667 7435 9673
rect 12250 9664 12256 9716
rect 12308 9704 12314 9716
rect 12437 9707 12495 9713
rect 12437 9704 12449 9707
rect 12308 9676 12449 9704
rect 12308 9664 12314 9676
rect 12437 9673 12449 9676
rect 12483 9673 12495 9707
rect 12437 9667 12495 9673
rect 12894 9664 12900 9716
rect 12952 9664 12958 9716
rect 8389 9639 8447 9645
rect 8389 9605 8401 9639
rect 8435 9605 8447 9639
rect 8389 9599 8447 9605
rect 7561 9503 7619 9509
rect 7561 9469 7573 9503
rect 7607 9500 7619 9503
rect 8404 9500 8432 9599
rect 8938 9528 8944 9580
rect 8996 9528 9002 9580
rect 12544 9540 13032 9568
rect 12544 9512 12572 9540
rect 7607 9472 8432 9500
rect 7607 9469 7619 9472
rect 7561 9463 7619 9469
rect 9030 9460 9036 9512
rect 9088 9500 9094 9512
rect 9401 9503 9459 9509
rect 9401 9500 9413 9503
rect 9088 9472 9413 9500
rect 9088 9460 9094 9472
rect 9401 9469 9413 9472
rect 9447 9469 9459 9503
rect 9401 9463 9459 9469
rect 9490 9460 9496 9512
rect 9548 9500 9554 9512
rect 9677 9503 9735 9509
rect 9677 9500 9689 9503
rect 9548 9472 9689 9500
rect 9548 9460 9554 9472
rect 9677 9469 9689 9472
rect 9723 9469 9735 9503
rect 9677 9463 9735 9469
rect 12345 9503 12403 9509
rect 12345 9469 12357 9503
rect 12391 9500 12403 9503
rect 12434 9500 12440 9512
rect 12391 9472 12440 9500
rect 12391 9469 12403 9472
rect 12345 9463 12403 9469
rect 12434 9460 12440 9472
rect 12492 9460 12498 9512
rect 12526 9460 12532 9512
rect 12584 9460 12590 9512
rect 12802 9460 12808 9512
rect 12860 9460 12866 9512
rect 13004 9509 13032 9540
rect 12989 9503 13047 9509
rect 12989 9469 13001 9503
rect 13035 9469 13047 9503
rect 12989 9463 13047 9469
rect 15010 9460 15016 9512
rect 15068 9460 15074 9512
rect 7006 9392 7012 9444
rect 7064 9432 7070 9444
rect 11425 9435 11483 9441
rect 11425 9432 11437 9435
rect 7064 9404 11437 9432
rect 7064 9392 7070 9404
rect 11425 9401 11437 9404
rect 11471 9432 11483 9435
rect 11471 9404 13032 9432
rect 11471 9401 11483 9404
rect 11425 9395 11483 9401
rect 13004 9376 13032 9404
rect 8754 9324 8760 9376
rect 8812 9324 8818 9376
rect 8846 9324 8852 9376
rect 8904 9324 8910 9376
rect 9493 9367 9551 9373
rect 9493 9333 9505 9367
rect 9539 9364 9551 9367
rect 9674 9364 9680 9376
rect 9539 9336 9680 9364
rect 9539 9333 9551 9336
rect 9493 9327 9551 9333
rect 9674 9324 9680 9336
rect 9732 9324 9738 9376
rect 12986 9324 12992 9376
rect 13044 9324 13050 9376
rect 552 9274 15520 9296
rect 552 9222 4100 9274
rect 4152 9222 4164 9274
rect 4216 9222 4228 9274
rect 4280 9222 4292 9274
rect 4344 9222 4356 9274
rect 4408 9222 7802 9274
rect 7854 9222 7866 9274
rect 7918 9222 7930 9274
rect 7982 9222 7994 9274
rect 8046 9222 8058 9274
rect 8110 9222 11504 9274
rect 11556 9222 11568 9274
rect 11620 9222 11632 9274
rect 11684 9222 11696 9274
rect 11748 9222 11760 9274
rect 11812 9222 15206 9274
rect 15258 9222 15270 9274
rect 15322 9222 15334 9274
rect 15386 9222 15398 9274
rect 15450 9222 15462 9274
rect 15514 9222 15520 9274
rect 552 9200 15520 9222
rect 8846 9120 8852 9172
rect 8904 9160 8910 9172
rect 8941 9163 8999 9169
rect 8941 9160 8953 9163
rect 8904 9132 8953 9160
rect 8904 9120 8910 9132
rect 8941 9129 8953 9132
rect 8987 9160 8999 9163
rect 12345 9163 12403 9169
rect 8987 9132 12296 9160
rect 8987 9129 8999 9132
rect 8941 9123 8999 9129
rect 8662 9092 8668 9104
rect 8050 9064 8668 9092
rect 8662 9052 8668 9064
rect 8720 9052 8726 9104
rect 10413 9095 10471 9101
rect 10413 9092 10425 9095
rect 9692 9064 10425 9092
rect 9692 9036 9720 9064
rect 10413 9061 10425 9064
rect 10459 9061 10471 9095
rect 10413 9055 10471 9061
rect 6641 9027 6699 9033
rect 6641 8993 6653 9027
rect 6687 9024 6699 9027
rect 6914 9024 6920 9036
rect 6687 8996 6920 9024
rect 6687 8993 6699 8996
rect 6641 8987 6699 8993
rect 6914 8984 6920 8996
rect 6972 8984 6978 9036
rect 7009 9027 7067 9033
rect 7009 8993 7021 9027
rect 7055 9024 7067 9027
rect 7098 9024 7104 9036
rect 7055 8996 7104 9024
rect 7055 8993 7067 8996
rect 7009 8987 7067 8993
rect 7098 8984 7104 8996
rect 7156 8984 7162 9036
rect 8754 8984 8760 9036
rect 8812 9024 8818 9036
rect 8812 8996 9444 9024
rect 8812 8984 8818 8996
rect 9416 8968 9444 8996
rect 9674 8984 9680 9036
rect 9732 8984 9738 9036
rect 9766 8984 9772 9036
rect 9824 8984 9830 9036
rect 10226 9033 10232 9036
rect 10219 9027 10232 9033
rect 10219 9024 10231 9027
rect 10187 8996 10231 9024
rect 10219 8993 10231 8996
rect 10219 8987 10232 8993
rect 10226 8984 10232 8987
rect 10284 8984 10290 9036
rect 10502 8984 10508 9036
rect 10560 9024 10566 9036
rect 11422 9024 11428 9036
rect 10560 8996 11428 9024
rect 10560 8984 10566 8996
rect 11422 8984 11428 8996
rect 11480 8984 11486 9036
rect 12158 8984 12164 9036
rect 12216 8984 12222 9036
rect 8435 8959 8493 8965
rect 8435 8925 8447 8959
rect 8481 8956 8493 8959
rect 9030 8956 9036 8968
rect 8481 8928 9036 8956
rect 8481 8925 8493 8928
rect 8435 8919 8493 8925
rect 9030 8916 9036 8928
rect 9088 8916 9094 8968
rect 9217 8959 9275 8965
rect 9217 8925 9229 8959
rect 9263 8956 9275 8959
rect 9306 8956 9312 8968
rect 9263 8928 9312 8956
rect 9263 8925 9275 8928
rect 9217 8919 9275 8925
rect 9306 8916 9312 8928
rect 9364 8916 9370 8968
rect 9398 8916 9404 8968
rect 9456 8956 9462 8968
rect 9784 8956 9812 8984
rect 9456 8928 9812 8956
rect 9456 8916 9462 8928
rect 10042 8916 10048 8968
rect 10100 8916 10106 8968
rect 10137 8959 10195 8965
rect 10137 8925 10149 8959
rect 10183 8925 10195 8959
rect 12268 8956 12296 9132
rect 12345 9129 12357 9163
rect 12391 9160 12403 9163
rect 12526 9160 12532 9172
rect 12391 9132 12532 9160
rect 12391 9129 12403 9132
rect 12345 9123 12403 9129
rect 12526 9120 12532 9132
rect 12584 9120 12590 9172
rect 13170 9052 13176 9104
rect 13228 9092 13234 9104
rect 13265 9095 13323 9101
rect 13265 9092 13277 9095
rect 13228 9064 13277 9092
rect 13228 9052 13234 9064
rect 13265 9061 13277 9064
rect 13311 9061 13323 9095
rect 13265 9055 13323 9061
rect 13722 9052 13728 9104
rect 13780 9052 13786 9104
rect 12342 8984 12348 9036
rect 12400 8984 12406 9036
rect 12986 8984 12992 9036
rect 13044 8984 13050 9036
rect 15013 8959 15071 8965
rect 15013 8956 15025 8959
rect 12268 8928 15025 8956
rect 10137 8919 10195 8925
rect 15013 8925 15025 8928
rect 15059 8956 15071 8959
rect 15562 8956 15568 8968
rect 15059 8928 15568 8956
rect 15059 8925 15071 8928
rect 15013 8919 15071 8925
rect 10152 8888 10180 8919
rect 15562 8916 15568 8928
rect 15620 8916 15626 8968
rect 10229 8891 10287 8897
rect 10229 8888 10241 8891
rect 10152 8860 10241 8888
rect 10229 8857 10241 8860
rect 10275 8857 10287 8891
rect 10229 8851 10287 8857
rect 8570 8780 8576 8832
rect 8628 8780 8634 8832
rect 9493 8823 9551 8829
rect 9493 8789 9505 8823
rect 9539 8820 9551 8823
rect 10686 8820 10692 8832
rect 9539 8792 10692 8820
rect 9539 8789 9551 8792
rect 9493 8783 9551 8789
rect 10686 8780 10692 8792
rect 10744 8780 10750 8832
rect 552 8730 15364 8752
rect 552 8678 2249 8730
rect 2301 8678 2313 8730
rect 2365 8678 2377 8730
rect 2429 8678 2441 8730
rect 2493 8678 2505 8730
rect 2557 8678 5951 8730
rect 6003 8678 6015 8730
rect 6067 8678 6079 8730
rect 6131 8678 6143 8730
rect 6195 8678 6207 8730
rect 6259 8678 9653 8730
rect 9705 8678 9717 8730
rect 9769 8678 9781 8730
rect 9833 8678 9845 8730
rect 9897 8678 9909 8730
rect 9961 8678 13355 8730
rect 13407 8678 13419 8730
rect 13471 8678 13483 8730
rect 13535 8678 13547 8730
rect 13599 8678 13611 8730
rect 13663 8678 15364 8730
rect 552 8656 15364 8678
rect 7098 8576 7104 8628
rect 7156 8576 7162 8628
rect 10226 8576 10232 8628
rect 10284 8616 10290 8628
rect 10870 8616 10876 8628
rect 10284 8588 10876 8616
rect 10284 8576 10290 8588
rect 10870 8576 10876 8588
rect 10928 8576 10934 8628
rect 11146 8576 11152 8628
rect 11204 8576 11210 8628
rect 9861 8551 9919 8557
rect 9861 8517 9873 8551
rect 9907 8517 9919 8551
rect 9861 8511 9919 8517
rect 10505 8551 10563 8557
rect 10505 8517 10517 8551
rect 10551 8548 10563 8551
rect 11793 8551 11851 8557
rect 10551 8520 11468 8548
rect 10551 8517 10563 8520
rect 10505 8511 10563 8517
rect 9398 8440 9404 8492
rect 9456 8440 9462 8492
rect 9876 8480 9904 8511
rect 9876 8452 10640 8480
rect 7285 8415 7343 8421
rect 7285 8381 7297 8415
rect 7331 8412 7343 8415
rect 8570 8412 8576 8424
rect 7331 8384 8576 8412
rect 7331 8381 7343 8384
rect 7285 8375 7343 8381
rect 8570 8372 8576 8384
rect 8628 8372 8634 8424
rect 9030 8372 9036 8424
rect 9088 8412 9094 8424
rect 9493 8415 9551 8421
rect 9493 8412 9505 8415
rect 9088 8384 9505 8412
rect 9088 8372 9094 8384
rect 9493 8381 9505 8384
rect 9539 8381 9551 8415
rect 9493 8375 9551 8381
rect 10226 8372 10232 8424
rect 10284 8372 10290 8424
rect 10502 8304 10508 8356
rect 10560 8304 10566 8356
rect 10612 8344 10640 8452
rect 10686 8440 10692 8492
rect 10744 8440 10750 8492
rect 10870 8440 10876 8492
rect 10928 8480 10934 8492
rect 11238 8480 11244 8492
rect 10928 8452 11244 8480
rect 10928 8440 10934 8452
rect 11238 8440 11244 8452
rect 11296 8440 11302 8492
rect 11333 8483 11391 8489
rect 11333 8449 11345 8483
rect 11379 8449 11391 8483
rect 11333 8443 11391 8449
rect 10778 8372 10784 8424
rect 10836 8372 10842 8424
rect 10965 8415 11023 8421
rect 10965 8381 10977 8415
rect 11011 8412 11023 8415
rect 11348 8412 11376 8443
rect 11440 8421 11468 8520
rect 11793 8517 11805 8551
rect 11839 8517 11851 8551
rect 11793 8511 11851 8517
rect 11808 8480 11836 8511
rect 12158 8480 12164 8492
rect 11808 8452 12164 8480
rect 12158 8440 12164 8452
rect 12216 8440 12222 8492
rect 11011 8384 11376 8412
rect 11425 8415 11483 8421
rect 11011 8381 11023 8384
rect 10965 8375 11023 8381
rect 11425 8381 11437 8415
rect 11471 8381 11483 8415
rect 11425 8375 11483 8381
rect 12253 8415 12311 8421
rect 12253 8381 12265 8415
rect 12299 8412 12311 8415
rect 12342 8412 12348 8424
rect 12299 8384 12348 8412
rect 12299 8381 12311 8384
rect 12253 8375 12311 8381
rect 10980 8344 11008 8375
rect 12342 8372 12348 8384
rect 12400 8372 12406 8424
rect 15013 8415 15071 8421
rect 15013 8381 15025 8415
rect 15059 8412 15071 8415
rect 15654 8412 15660 8424
rect 15059 8384 15660 8412
rect 15059 8381 15071 8384
rect 15013 8375 15071 8381
rect 15654 8372 15660 8384
rect 15712 8372 15718 8424
rect 10612 8316 11008 8344
rect 10321 8279 10379 8285
rect 10321 8245 10333 8279
rect 10367 8276 10379 8279
rect 10778 8276 10784 8288
rect 10367 8248 10784 8276
rect 10367 8245 10379 8248
rect 10321 8239 10379 8245
rect 10778 8236 10784 8248
rect 10836 8236 10842 8288
rect 12618 8236 12624 8288
rect 12676 8236 12682 8288
rect 552 8186 15520 8208
rect 552 8134 4100 8186
rect 4152 8134 4164 8186
rect 4216 8134 4228 8186
rect 4280 8134 4292 8186
rect 4344 8134 4356 8186
rect 4408 8134 7802 8186
rect 7854 8134 7866 8186
rect 7918 8134 7930 8186
rect 7982 8134 7994 8186
rect 8046 8134 8058 8186
rect 8110 8134 11504 8186
rect 11556 8134 11568 8186
rect 11620 8134 11632 8186
rect 11684 8134 11696 8186
rect 11748 8134 11760 8186
rect 11812 8134 15206 8186
rect 15258 8134 15270 8186
rect 15322 8134 15334 8186
rect 15386 8134 15398 8186
rect 15450 8134 15462 8186
rect 15514 8134 15520 8186
rect 552 8112 15520 8134
rect 8757 8075 8815 8081
rect 8757 8041 8769 8075
rect 8803 8072 8815 8075
rect 8803 8044 9352 8072
rect 8803 8041 8815 8044
rect 8757 8035 8815 8041
rect 8662 8004 8668 8016
rect 8510 7976 8668 8004
rect 8662 7964 8668 7976
rect 8720 8004 8726 8016
rect 9214 8004 9220 8016
rect 8720 7976 9220 8004
rect 8720 7964 8726 7976
rect 9214 7964 9220 7976
rect 9272 7964 9278 8016
rect 7006 7896 7012 7948
rect 7064 7896 7070 7948
rect 9324 7945 9352 8044
rect 10502 8032 10508 8084
rect 10560 8072 10566 8084
rect 10781 8075 10839 8081
rect 10781 8072 10793 8075
rect 10560 8044 10793 8072
rect 10560 8032 10566 8044
rect 10781 8041 10793 8044
rect 10827 8041 10839 8075
rect 10781 8035 10839 8041
rect 9309 7939 9367 7945
rect 9309 7905 9321 7939
rect 9355 7936 9367 7939
rect 10796 7936 10824 8035
rect 10870 8032 10876 8084
rect 10928 8072 10934 8084
rect 11609 8075 11667 8081
rect 11609 8072 11621 8075
rect 10928 8044 11621 8072
rect 10928 8032 10934 8044
rect 11609 8041 11621 8044
rect 11655 8041 11667 8075
rect 11609 8035 11667 8041
rect 13170 8004 13176 8016
rect 12544 7976 13176 8004
rect 12544 7945 12572 7976
rect 13170 7964 13176 7976
rect 13228 7964 13234 8016
rect 13722 7964 13728 8016
rect 13780 7964 13786 8016
rect 15010 7964 15016 8016
rect 15068 7964 15074 8016
rect 11517 7939 11575 7945
rect 11517 7936 11529 7939
rect 9355 7908 9628 7936
rect 10796 7908 11529 7936
rect 9355 7905 9367 7908
rect 9309 7899 9367 7905
rect 7282 7828 7288 7880
rect 7340 7828 7346 7880
rect 8938 7828 8944 7880
rect 8996 7828 9002 7880
rect 9214 7828 9220 7880
rect 9272 7868 9278 7880
rect 9401 7871 9459 7877
rect 9401 7868 9413 7871
rect 9272 7840 9413 7868
rect 9272 7828 9278 7840
rect 9401 7837 9413 7840
rect 9447 7837 9459 7871
rect 9401 7831 9459 7837
rect 9493 7871 9551 7877
rect 9493 7837 9505 7871
rect 9539 7837 9551 7871
rect 9600 7868 9628 7908
rect 11517 7905 11529 7908
rect 11563 7905 11575 7939
rect 11517 7899 11575 7905
rect 11701 7939 11759 7945
rect 11701 7905 11713 7939
rect 11747 7905 11759 7939
rect 11701 7899 11759 7905
rect 12529 7939 12587 7945
rect 12529 7905 12541 7939
rect 12575 7905 12587 7939
rect 12529 7899 12587 7905
rect 10318 7868 10324 7880
rect 9600 7840 10324 7868
rect 9493 7831 9551 7837
rect 8956 7800 8984 7828
rect 9508 7800 9536 7831
rect 10318 7828 10324 7840
rect 10376 7828 10382 7880
rect 10965 7871 11023 7877
rect 10965 7837 10977 7871
rect 11011 7837 11023 7871
rect 10965 7831 11023 7837
rect 11425 7871 11483 7877
rect 11425 7837 11437 7871
rect 11471 7868 11483 7871
rect 11716 7868 11744 7899
rect 12986 7896 12992 7948
rect 13044 7896 13050 7948
rect 11471 7840 11744 7868
rect 11471 7837 11483 7840
rect 11425 7831 11483 7837
rect 8956 7772 9536 7800
rect 10042 7760 10048 7812
rect 10100 7800 10106 7812
rect 10594 7800 10600 7812
rect 10100 7772 10600 7800
rect 10100 7760 10106 7772
rect 10594 7760 10600 7772
rect 10652 7800 10658 7812
rect 10980 7800 11008 7831
rect 12618 7828 12624 7880
rect 12676 7828 12682 7880
rect 12897 7871 12955 7877
rect 12897 7837 12909 7871
rect 12943 7868 12955 7871
rect 13265 7871 13323 7877
rect 13265 7868 13277 7871
rect 12943 7840 13277 7868
rect 12943 7837 12955 7840
rect 12897 7831 12955 7837
rect 13265 7837 13277 7840
rect 13311 7837 13323 7871
rect 13265 7831 13323 7837
rect 10652 7772 11008 7800
rect 11333 7803 11391 7809
rect 10652 7760 10658 7772
rect 11333 7769 11345 7803
rect 11379 7800 11391 7803
rect 12342 7800 12348 7812
rect 11379 7772 12348 7800
rect 11379 7769 11391 7772
rect 11333 7763 11391 7769
rect 8938 7692 8944 7744
rect 8996 7692 9002 7744
rect 10318 7692 10324 7744
rect 10376 7732 10382 7744
rect 11348 7732 11376 7763
rect 12342 7760 12348 7772
rect 12400 7760 12406 7812
rect 10376 7704 11376 7732
rect 10376 7692 10382 7704
rect 552 7642 15364 7664
rect 552 7590 2249 7642
rect 2301 7590 2313 7642
rect 2365 7590 2377 7642
rect 2429 7590 2441 7642
rect 2493 7590 2505 7642
rect 2557 7590 5951 7642
rect 6003 7590 6015 7642
rect 6067 7590 6079 7642
rect 6131 7590 6143 7642
rect 6195 7590 6207 7642
rect 6259 7590 9653 7642
rect 9705 7590 9717 7642
rect 9769 7590 9781 7642
rect 9833 7590 9845 7642
rect 9897 7590 9909 7642
rect 9961 7590 13355 7642
rect 13407 7590 13419 7642
rect 13471 7590 13483 7642
rect 13535 7590 13547 7642
rect 13599 7590 13611 7642
rect 13663 7590 15364 7642
rect 552 7568 15364 7590
rect 7282 7488 7288 7540
rect 7340 7528 7346 7540
rect 7469 7531 7527 7537
rect 7469 7528 7481 7531
rect 7340 7500 7481 7528
rect 7340 7488 7346 7500
rect 7469 7497 7481 7500
rect 7515 7497 7527 7531
rect 7469 7491 7527 7497
rect 12621 7531 12679 7537
rect 12621 7497 12633 7531
rect 12667 7528 12679 7531
rect 12802 7528 12808 7540
rect 12667 7500 12808 7528
rect 12667 7497 12679 7500
rect 12621 7491 12679 7497
rect 12802 7488 12808 7500
rect 12860 7488 12866 7540
rect 13170 7488 13176 7540
rect 13228 7528 13234 7540
rect 13541 7531 13599 7537
rect 13541 7528 13553 7531
rect 13228 7500 13553 7528
rect 13228 7488 13234 7500
rect 13541 7497 13553 7500
rect 13587 7497 13599 7531
rect 13541 7491 13599 7497
rect 13262 7460 13268 7472
rect 11532 7432 13268 7460
rect 7653 7327 7711 7333
rect 7653 7293 7665 7327
rect 7699 7324 7711 7327
rect 8938 7324 8944 7336
rect 7699 7296 8944 7324
rect 7699 7293 7711 7296
rect 7653 7287 7711 7293
rect 8938 7284 8944 7296
rect 8996 7284 9002 7336
rect 9306 7284 9312 7336
rect 9364 7284 9370 7336
rect 11532 7333 11560 7432
rect 13262 7420 13268 7432
rect 13320 7420 13326 7472
rect 12618 7352 12624 7404
rect 12676 7392 12682 7404
rect 14001 7395 14059 7401
rect 14001 7392 14013 7395
rect 12676 7364 13216 7392
rect 12676 7352 12682 7364
rect 11517 7327 11575 7333
rect 11517 7293 11529 7327
rect 11563 7293 11575 7327
rect 11517 7287 11575 7293
rect 12802 7284 12808 7336
rect 12860 7324 12866 7336
rect 13188 7333 13216 7364
rect 13280 7364 14013 7392
rect 13280 7336 13308 7364
rect 14001 7361 14013 7364
rect 14047 7361 14059 7395
rect 14001 7355 14059 7361
rect 13173 7327 13231 7333
rect 12860 7296 13124 7324
rect 12860 7284 12866 7296
rect 9582 7216 9588 7268
rect 9640 7256 9646 7268
rect 9769 7259 9827 7265
rect 9769 7256 9781 7259
rect 9640 7228 9781 7256
rect 9640 7216 9646 7228
rect 9769 7225 9781 7228
rect 9815 7225 9827 7259
rect 9769 7219 9827 7225
rect 12894 7216 12900 7268
rect 12952 7216 12958 7268
rect 12989 7259 13047 7265
rect 12989 7225 13001 7259
rect 13035 7225 13047 7259
rect 13096 7256 13124 7296
rect 13173 7293 13185 7327
rect 13219 7293 13231 7327
rect 13173 7287 13231 7293
rect 13262 7284 13268 7336
rect 13320 7284 13326 7336
rect 13725 7327 13783 7333
rect 13725 7293 13737 7327
rect 13771 7293 13783 7327
rect 13725 7287 13783 7293
rect 13740 7256 13768 7287
rect 13814 7284 13820 7336
rect 13872 7284 13878 7336
rect 13909 7327 13967 7333
rect 13909 7293 13921 7327
rect 13955 7293 13967 7327
rect 13909 7287 13967 7293
rect 13096 7228 13768 7256
rect 12989 7219 13047 7225
rect 9122 7148 9128 7200
rect 9180 7148 9186 7200
rect 13004 7188 13032 7219
rect 13722 7188 13728 7200
rect 13004 7160 13728 7188
rect 13722 7148 13728 7160
rect 13780 7188 13786 7200
rect 13924 7188 13952 7287
rect 13780 7160 13952 7188
rect 13780 7148 13786 7160
rect 552 7098 15520 7120
rect 552 7046 4100 7098
rect 4152 7046 4164 7098
rect 4216 7046 4228 7098
rect 4280 7046 4292 7098
rect 4344 7046 4356 7098
rect 4408 7046 7802 7098
rect 7854 7046 7866 7098
rect 7918 7046 7930 7098
rect 7982 7046 7994 7098
rect 8046 7046 8058 7098
rect 8110 7046 11504 7098
rect 11556 7046 11568 7098
rect 11620 7046 11632 7098
rect 11684 7046 11696 7098
rect 11748 7046 11760 7098
rect 11812 7046 15206 7098
rect 15258 7046 15270 7098
rect 15322 7046 15334 7098
rect 15386 7046 15398 7098
rect 15450 7046 15462 7098
rect 15514 7046 15520 7098
rect 552 7024 15520 7046
rect 10594 6993 10600 6996
rect 10551 6987 10600 6993
rect 8220 6956 9444 6984
rect 8110 6916 8116 6928
rect 8050 6888 8116 6916
rect 8110 6876 8116 6888
rect 8168 6916 8174 6928
rect 8220 6916 8248 6956
rect 8168 6888 8248 6916
rect 9416 6916 9444 6956
rect 10551 6953 10563 6987
rect 10597 6953 10600 6987
rect 10551 6947 10600 6953
rect 10594 6944 10600 6947
rect 10652 6944 10658 6996
rect 12345 6919 12403 6925
rect 9416 6888 9522 6916
rect 8168 6876 8174 6888
rect 12345 6885 12357 6919
rect 12391 6916 12403 6919
rect 12391 6888 12848 6916
rect 12391 6885 12403 6888
rect 12345 6879 12403 6885
rect 12820 6860 12848 6888
rect 9122 6808 9128 6860
rect 9180 6808 9186 6860
rect 10870 6808 10876 6860
rect 10928 6848 10934 6860
rect 11149 6851 11207 6857
rect 11149 6848 11161 6851
rect 10928 6820 11161 6848
rect 10928 6808 10934 6820
rect 11149 6817 11161 6820
rect 11195 6817 11207 6851
rect 11149 6811 11207 6817
rect 11974 6808 11980 6860
rect 12032 6808 12038 6860
rect 12161 6851 12219 6857
rect 12161 6817 12173 6851
rect 12207 6848 12219 6851
rect 12253 6851 12311 6857
rect 12253 6848 12265 6851
rect 12207 6820 12265 6848
rect 12207 6817 12219 6820
rect 12161 6811 12219 6817
rect 12253 6817 12265 6820
rect 12299 6817 12311 6851
rect 12253 6811 12311 6817
rect 12437 6851 12495 6857
rect 12437 6817 12449 6851
rect 12483 6817 12495 6851
rect 12437 6811 12495 6817
rect 6546 6740 6552 6792
rect 6604 6740 6610 6792
rect 6822 6740 6828 6792
rect 6880 6740 6886 6792
rect 8754 6740 8760 6792
rect 8812 6740 8818 6792
rect 11238 6740 11244 6792
rect 11296 6740 11302 6792
rect 11517 6783 11575 6789
rect 11517 6749 11529 6783
rect 11563 6780 11575 6783
rect 12176 6780 12204 6811
rect 11563 6752 12204 6780
rect 11563 6749 11575 6752
rect 11517 6743 11575 6749
rect 11974 6672 11980 6724
rect 12032 6712 12038 6724
rect 12452 6712 12480 6811
rect 12802 6808 12808 6860
rect 12860 6848 12866 6860
rect 12897 6851 12955 6857
rect 12897 6848 12909 6851
rect 12860 6820 12909 6848
rect 12860 6808 12866 6820
rect 12897 6817 12909 6820
rect 12943 6817 12955 6851
rect 12897 6811 12955 6817
rect 12032 6684 12480 6712
rect 12032 6672 12038 6684
rect 8294 6604 8300 6656
rect 8352 6604 8358 6656
rect 12161 6647 12219 6653
rect 12161 6613 12173 6647
rect 12207 6644 12219 6647
rect 13173 6647 13231 6653
rect 13173 6644 13185 6647
rect 12207 6616 13185 6644
rect 12207 6613 12219 6616
rect 12161 6607 12219 6613
rect 13173 6613 13185 6616
rect 13219 6644 13231 6647
rect 13262 6644 13268 6656
rect 13219 6616 13268 6644
rect 13219 6613 13231 6616
rect 13173 6607 13231 6613
rect 13262 6604 13268 6616
rect 13320 6604 13326 6656
rect 13357 6647 13415 6653
rect 13357 6613 13369 6647
rect 13403 6644 13415 6647
rect 13906 6644 13912 6656
rect 13403 6616 13912 6644
rect 13403 6613 13415 6616
rect 13357 6607 13415 6613
rect 13906 6604 13912 6616
rect 13964 6604 13970 6656
rect 552 6554 15364 6576
rect 552 6502 2249 6554
rect 2301 6502 2313 6554
rect 2365 6502 2377 6554
rect 2429 6502 2441 6554
rect 2493 6502 2505 6554
rect 2557 6502 5951 6554
rect 6003 6502 6015 6554
rect 6067 6502 6079 6554
rect 6131 6502 6143 6554
rect 6195 6502 6207 6554
rect 6259 6502 9653 6554
rect 9705 6502 9717 6554
rect 9769 6502 9781 6554
rect 9833 6502 9845 6554
rect 9897 6502 9909 6554
rect 9961 6502 13355 6554
rect 13407 6502 13419 6554
rect 13471 6502 13483 6554
rect 13535 6502 13547 6554
rect 13599 6502 13611 6554
rect 13663 6502 15364 6554
rect 552 6480 15364 6502
rect 6822 6400 6828 6452
rect 6880 6440 6886 6452
rect 7101 6443 7159 6449
rect 7101 6440 7113 6443
rect 6880 6412 7113 6440
rect 6880 6400 6886 6412
rect 7101 6409 7113 6412
rect 7147 6409 7159 6443
rect 7101 6403 7159 6409
rect 8021 6443 8079 6449
rect 8021 6409 8033 6443
rect 8067 6440 8079 6443
rect 8110 6440 8116 6452
rect 8067 6412 8116 6440
rect 8067 6409 8079 6412
rect 8021 6403 8079 6409
rect 8110 6400 8116 6412
rect 8168 6400 8174 6452
rect 9306 6400 9312 6452
rect 9364 6400 9370 6452
rect 8389 6375 8447 6381
rect 8389 6341 8401 6375
rect 8435 6341 8447 6375
rect 8389 6335 8447 6341
rect 7285 6239 7343 6245
rect 7285 6205 7297 6239
rect 7331 6236 7343 6239
rect 8404 6236 8432 6335
rect 9030 6264 9036 6316
rect 9088 6264 9094 6316
rect 9398 6264 9404 6316
rect 9456 6304 9462 6316
rect 9861 6307 9919 6313
rect 9861 6304 9873 6307
rect 9456 6276 9873 6304
rect 9456 6264 9462 6276
rect 9861 6273 9873 6276
rect 9907 6273 9919 6307
rect 9861 6267 9919 6273
rect 13265 6307 13323 6313
rect 13265 6273 13277 6307
rect 13311 6304 13323 6307
rect 13817 6307 13875 6313
rect 13817 6304 13829 6307
rect 13311 6276 13829 6304
rect 13311 6273 13323 6276
rect 13265 6267 13323 6273
rect 13817 6273 13829 6276
rect 13863 6273 13875 6307
rect 13817 6267 13875 6273
rect 7331 6208 8432 6236
rect 7331 6205 7343 6208
rect 7285 6199 7343 6205
rect 9214 6196 9220 6248
rect 9272 6236 9278 6248
rect 9677 6239 9735 6245
rect 9677 6236 9689 6239
rect 9272 6208 9689 6236
rect 9272 6196 9278 6208
rect 9677 6205 9689 6208
rect 9723 6205 9735 6239
rect 9677 6199 9735 6205
rect 9769 6239 9827 6245
rect 9769 6205 9781 6239
rect 9815 6236 9827 6239
rect 10594 6236 10600 6248
rect 9815 6208 10600 6236
rect 9815 6205 9827 6208
rect 9769 6199 9827 6205
rect 10594 6196 10600 6208
rect 10652 6196 10658 6248
rect 12894 6196 12900 6248
rect 12952 6236 12958 6248
rect 13173 6239 13231 6245
rect 13173 6236 13185 6239
rect 12952 6208 13185 6236
rect 12952 6196 12958 6208
rect 13173 6205 13185 6208
rect 13219 6205 13231 6239
rect 13173 6199 13231 6205
rect 13357 6239 13415 6245
rect 13357 6205 13369 6239
rect 13403 6236 13415 6239
rect 13722 6236 13728 6248
rect 13403 6208 13728 6236
rect 13403 6205 13415 6208
rect 13357 6199 13415 6205
rect 8113 6171 8171 6177
rect 8113 6137 8125 6171
rect 8159 6137 8171 6171
rect 8113 6131 8171 6137
rect 8128 6100 8156 6131
rect 8294 6128 8300 6180
rect 8352 6168 8358 6180
rect 8757 6171 8815 6177
rect 8757 6168 8769 6171
rect 8352 6140 8769 6168
rect 8352 6128 8358 6140
rect 8757 6137 8769 6140
rect 8803 6168 8815 6171
rect 9582 6168 9588 6180
rect 8803 6140 9588 6168
rect 8803 6137 8815 6140
rect 8757 6131 8815 6137
rect 9582 6128 9588 6140
rect 9640 6128 9646 6180
rect 13188 6168 13216 6199
rect 13722 6196 13728 6208
rect 13780 6196 13786 6248
rect 13906 6196 13912 6248
rect 13964 6196 13970 6248
rect 13814 6168 13820 6180
rect 13188 6140 13820 6168
rect 13814 6128 13820 6140
rect 13872 6128 13878 6180
rect 8386 6100 8392 6112
rect 8128 6072 8392 6100
rect 8386 6060 8392 6072
rect 8444 6060 8450 6112
rect 8849 6103 8907 6109
rect 8849 6069 8861 6103
rect 8895 6100 8907 6103
rect 9122 6100 9128 6112
rect 8895 6072 9128 6100
rect 8895 6069 8907 6072
rect 8849 6063 8907 6069
rect 9122 6060 9128 6072
rect 9180 6060 9186 6112
rect 13538 6060 13544 6112
rect 13596 6060 13602 6112
rect 552 6010 15520 6032
rect 552 5958 4100 6010
rect 4152 5958 4164 6010
rect 4216 5958 4228 6010
rect 4280 5958 4292 6010
rect 4344 5958 4356 6010
rect 4408 5958 7802 6010
rect 7854 5958 7866 6010
rect 7918 5958 7930 6010
rect 7982 5958 7994 6010
rect 8046 5958 8058 6010
rect 8110 5958 11504 6010
rect 11556 5958 11568 6010
rect 11620 5958 11632 6010
rect 11684 5958 11696 6010
rect 11748 5958 11760 6010
rect 11812 5958 15206 6010
rect 15258 5958 15270 6010
rect 15322 5958 15334 6010
rect 15386 5958 15398 6010
rect 15450 5958 15462 6010
rect 15514 5958 15520 6010
rect 552 5936 15520 5958
rect 9122 5856 9128 5908
rect 9180 5896 9186 5908
rect 15010 5896 15016 5908
rect 9180 5868 15016 5896
rect 9180 5856 9186 5868
rect 15010 5856 15016 5868
rect 15068 5856 15074 5908
rect 8202 5788 8208 5840
rect 8260 5788 8266 5840
rect 8619 5831 8677 5837
rect 8619 5797 8631 5831
rect 8665 5828 8677 5831
rect 9217 5831 9275 5837
rect 9217 5828 9229 5831
rect 8665 5800 9229 5828
rect 8665 5797 8677 5800
rect 8619 5791 8677 5797
rect 9217 5797 9229 5800
rect 9263 5797 9275 5831
rect 9217 5791 9275 5797
rect 13265 5831 13323 5837
rect 13265 5797 13277 5831
rect 13311 5828 13323 5831
rect 13538 5828 13544 5840
rect 13311 5800 13544 5828
rect 13311 5797 13323 5800
rect 13265 5791 13323 5797
rect 6546 5720 6552 5772
rect 6604 5760 6610 5772
rect 6825 5763 6883 5769
rect 6825 5760 6837 5763
rect 6604 5732 6837 5760
rect 6604 5720 6610 5732
rect 6825 5729 6837 5732
rect 6871 5760 6883 5763
rect 6871 5732 7328 5760
rect 6871 5729 6883 5732
rect 6825 5723 6883 5729
rect 7190 5652 7196 5704
rect 7248 5652 7254 5704
rect 7300 5692 7328 5732
rect 8754 5692 8760 5704
rect 7300 5664 8760 5692
rect 8754 5652 8760 5664
rect 8812 5652 8818 5704
rect 9232 5624 9260 5791
rect 13538 5788 13544 5800
rect 13596 5788 13602 5840
rect 13906 5788 13912 5840
rect 13964 5788 13970 5840
rect 9582 5720 9588 5772
rect 9640 5760 9646 5772
rect 9640 5732 10548 5760
rect 9640 5720 9646 5732
rect 9398 5652 9404 5704
rect 9456 5652 9462 5704
rect 10137 5695 10195 5701
rect 10137 5661 10149 5695
rect 10183 5661 10195 5695
rect 10137 5655 10195 5661
rect 9861 5627 9919 5633
rect 9861 5624 9873 5627
rect 9232 5596 9873 5624
rect 9861 5593 9873 5596
rect 9907 5624 9919 5627
rect 10152 5624 10180 5655
rect 10520 5633 10548 5732
rect 12986 5652 12992 5704
rect 13044 5652 13050 5704
rect 15010 5652 15016 5704
rect 15068 5652 15074 5704
rect 9907 5596 10180 5624
rect 10505 5627 10563 5633
rect 9907 5593 9919 5596
rect 9861 5587 9919 5593
rect 10505 5593 10517 5627
rect 10551 5624 10563 5627
rect 11974 5624 11980 5636
rect 10551 5596 11980 5624
rect 10551 5593 10563 5596
rect 10505 5587 10563 5593
rect 11974 5584 11980 5596
rect 12032 5584 12038 5636
rect 8757 5559 8815 5565
rect 8757 5525 8769 5559
rect 8803 5556 8815 5559
rect 8846 5556 8852 5568
rect 8803 5528 8852 5556
rect 8803 5525 8815 5528
rect 8757 5519 8815 5525
rect 8846 5516 8852 5528
rect 8904 5516 8910 5568
rect 10042 5516 10048 5568
rect 10100 5516 10106 5568
rect 10226 5516 10232 5568
rect 10284 5556 10290 5568
rect 10597 5559 10655 5565
rect 10597 5556 10609 5559
rect 10284 5528 10609 5556
rect 10284 5516 10290 5528
rect 10597 5525 10609 5528
rect 10643 5525 10655 5559
rect 10597 5519 10655 5525
rect 552 5466 15364 5488
rect 552 5414 2249 5466
rect 2301 5414 2313 5466
rect 2365 5414 2377 5466
rect 2429 5414 2441 5466
rect 2493 5414 2505 5466
rect 2557 5414 5951 5466
rect 6003 5414 6015 5466
rect 6067 5414 6079 5466
rect 6131 5414 6143 5466
rect 6195 5414 6207 5466
rect 6259 5414 9653 5466
rect 9705 5414 9717 5466
rect 9769 5414 9781 5466
rect 9833 5414 9845 5466
rect 9897 5414 9909 5466
rect 9961 5414 13355 5466
rect 13407 5414 13419 5466
rect 13471 5414 13483 5466
rect 13535 5414 13547 5466
rect 13599 5414 13611 5466
rect 13663 5414 15364 5466
rect 552 5392 15364 5414
rect 7190 5312 7196 5364
rect 7248 5352 7254 5364
rect 7285 5355 7343 5361
rect 7285 5352 7297 5355
rect 7248 5324 7297 5352
rect 7248 5312 7254 5324
rect 7285 5321 7297 5324
rect 7331 5321 7343 5355
rect 7285 5315 7343 5321
rect 11238 5312 11244 5364
rect 11296 5352 11302 5364
rect 11885 5355 11943 5361
rect 11885 5352 11897 5355
rect 11296 5324 11897 5352
rect 11296 5312 11302 5324
rect 11885 5321 11897 5324
rect 11931 5321 11943 5355
rect 11885 5315 11943 5321
rect 13633 5355 13691 5361
rect 13633 5321 13645 5355
rect 13679 5352 13691 5355
rect 13722 5352 13728 5364
rect 13679 5324 13728 5352
rect 13679 5321 13691 5324
rect 13633 5315 13691 5321
rect 13722 5312 13728 5324
rect 13780 5312 13786 5364
rect 8754 5244 8760 5296
rect 8812 5284 8818 5296
rect 12986 5284 12992 5296
rect 8812 5256 12992 5284
rect 8812 5244 8818 5256
rect 11164 5225 11192 5256
rect 12986 5244 12992 5256
rect 13044 5244 13050 5296
rect 11149 5219 11207 5225
rect 11149 5185 11161 5219
rect 11195 5185 11207 5219
rect 11149 5179 11207 5185
rect 12069 5219 12127 5225
rect 12069 5185 12081 5219
rect 12115 5185 12127 5219
rect 12713 5219 12771 5225
rect 12713 5216 12725 5219
rect 12069 5179 12127 5185
rect 12544 5188 12725 5216
rect 7469 5151 7527 5157
rect 7469 5117 7481 5151
rect 7515 5148 7527 5151
rect 8846 5148 8852 5160
rect 7515 5120 8852 5148
rect 7515 5117 7527 5120
rect 7469 5111 7527 5117
rect 8846 5108 8852 5120
rect 8904 5108 8910 5160
rect 9401 5151 9459 5157
rect 9401 5117 9413 5151
rect 9447 5148 9459 5151
rect 9490 5148 9496 5160
rect 9447 5120 9496 5148
rect 9447 5117 9459 5120
rect 9401 5111 9459 5117
rect 9490 5108 9496 5120
rect 9548 5108 9554 5160
rect 10042 5108 10048 5160
rect 10100 5148 10106 5160
rect 11241 5151 11299 5157
rect 11241 5148 11253 5151
rect 10100 5120 11253 5148
rect 10100 5108 10106 5120
rect 11241 5117 11253 5120
rect 11287 5117 11299 5151
rect 11241 5111 11299 5117
rect 11330 5108 11336 5160
rect 11388 5108 11394 5160
rect 11422 5108 11428 5160
rect 11480 5148 11486 5160
rect 11609 5151 11667 5157
rect 11609 5148 11621 5151
rect 11480 5120 11621 5148
rect 11480 5108 11486 5120
rect 11609 5117 11621 5120
rect 11655 5117 11667 5151
rect 11609 5111 11667 5117
rect 11701 5151 11759 5157
rect 11701 5117 11713 5151
rect 11747 5148 11759 5151
rect 12084 5148 12112 5179
rect 11747 5120 12112 5148
rect 11747 5117 11759 5120
rect 11701 5111 11759 5117
rect 11054 5040 11060 5092
rect 11112 5080 11118 5092
rect 11517 5083 11575 5089
rect 11517 5080 11529 5083
rect 11112 5052 11529 5080
rect 11112 5040 11118 5052
rect 11517 5049 11529 5052
rect 11563 5049 11575 5083
rect 11517 5043 11575 5049
rect 10686 4972 10692 5024
rect 10744 5012 10750 5024
rect 11716 5012 11744 5111
rect 12158 5108 12164 5160
rect 12216 5108 12222 5160
rect 12544 5021 12572 5188
rect 12713 5185 12725 5188
rect 12759 5216 12771 5219
rect 12759 5188 13584 5216
rect 12759 5185 12771 5188
rect 12713 5179 12771 5185
rect 12802 5108 12808 5160
rect 12860 5108 12866 5160
rect 13556 5157 13584 5188
rect 13541 5151 13599 5157
rect 13541 5117 13553 5151
rect 13587 5117 13599 5151
rect 13541 5111 13599 5117
rect 13722 5108 13728 5160
rect 13780 5108 13786 5160
rect 10744 4984 11744 5012
rect 12529 5015 12587 5021
rect 10744 4972 10750 4984
rect 12529 4981 12541 5015
rect 12575 4981 12587 5015
rect 12529 4975 12587 4981
rect 13170 4972 13176 5024
rect 13228 4972 13234 5024
rect 552 4922 15520 4944
rect 552 4870 4100 4922
rect 4152 4870 4164 4922
rect 4216 4870 4228 4922
rect 4280 4870 4292 4922
rect 4344 4870 4356 4922
rect 4408 4870 7802 4922
rect 7854 4870 7866 4922
rect 7918 4870 7930 4922
rect 7982 4870 7994 4922
rect 8046 4870 8058 4922
rect 8110 4870 11504 4922
rect 11556 4870 11568 4922
rect 11620 4870 11632 4922
rect 11684 4870 11696 4922
rect 11748 4870 11760 4922
rect 11812 4870 15206 4922
rect 15258 4870 15270 4922
rect 15322 4870 15334 4922
rect 15386 4870 15398 4922
rect 15450 4870 15462 4922
rect 15514 4870 15520 4922
rect 552 4848 15520 4870
rect 10045 4811 10103 4817
rect 10045 4777 10057 4811
rect 10091 4808 10103 4811
rect 10686 4808 10692 4820
rect 10091 4780 10692 4808
rect 10091 4777 10103 4780
rect 10045 4771 10103 4777
rect 10686 4768 10692 4780
rect 10744 4768 10750 4820
rect 10781 4811 10839 4817
rect 10781 4777 10793 4811
rect 10827 4808 10839 4811
rect 11330 4808 11336 4820
rect 10827 4780 11336 4808
rect 10827 4777 10839 4780
rect 10781 4771 10839 4777
rect 11330 4768 11336 4780
rect 11388 4768 11394 4820
rect 10597 4743 10655 4749
rect 10597 4709 10609 4743
rect 10643 4740 10655 4743
rect 12345 4743 12403 4749
rect 12345 4740 12357 4743
rect 10643 4712 12357 4740
rect 10643 4709 10655 4712
rect 10597 4703 10655 4709
rect 12345 4709 12357 4712
rect 12391 4740 12403 4743
rect 12802 4740 12808 4752
rect 12391 4712 12808 4740
rect 12391 4709 12403 4712
rect 12345 4703 12403 4709
rect 12802 4700 12808 4712
rect 12860 4700 12866 4752
rect 9214 4632 9220 4684
rect 9272 4632 9278 4684
rect 9953 4675 10011 4681
rect 9953 4641 9965 4675
rect 9999 4672 10011 4675
rect 10042 4672 10048 4684
rect 9999 4644 10048 4672
rect 9999 4641 10011 4644
rect 9953 4635 10011 4641
rect 10042 4632 10048 4644
rect 10100 4632 10106 4684
rect 10137 4675 10195 4681
rect 10137 4641 10149 4675
rect 10183 4672 10195 4675
rect 10226 4672 10232 4684
rect 10183 4644 10232 4672
rect 10183 4641 10195 4644
rect 10137 4635 10195 4641
rect 10226 4632 10232 4644
rect 10284 4632 10290 4684
rect 11149 4675 11207 4681
rect 11149 4641 11161 4675
rect 11195 4672 11207 4675
rect 11238 4672 11244 4684
rect 11195 4644 11244 4672
rect 11195 4641 11207 4644
rect 11149 4635 11207 4641
rect 11238 4632 11244 4644
rect 11296 4632 11302 4684
rect 11330 4632 11336 4684
rect 11388 4632 11394 4684
rect 11422 4632 11428 4684
rect 11480 4632 11486 4684
rect 11514 4632 11520 4684
rect 11572 4672 11578 4684
rect 12437 4675 12495 4681
rect 12437 4672 12449 4675
rect 11572 4644 12449 4672
rect 11572 4632 11578 4644
rect 12437 4641 12449 4644
rect 12483 4672 12495 4675
rect 13722 4672 13728 4684
rect 12483 4644 13728 4672
rect 12483 4641 12495 4644
rect 12437 4635 12495 4641
rect 13722 4632 13728 4644
rect 13780 4632 13786 4684
rect 13906 4632 13912 4684
rect 13964 4632 13970 4684
rect 11054 4564 11060 4616
rect 11112 4604 11118 4616
rect 11348 4604 11376 4632
rect 11112 4576 11376 4604
rect 11112 4564 11118 4576
rect 11149 4539 11207 4545
rect 11149 4505 11161 4539
rect 11195 4536 11207 4539
rect 12158 4536 12164 4548
rect 11195 4508 12164 4536
rect 11195 4505 11207 4508
rect 11149 4499 11207 4505
rect 12158 4496 12164 4508
rect 12216 4496 12222 4548
rect 8938 4428 8944 4480
rect 8996 4468 9002 4480
rect 9033 4471 9091 4477
rect 9033 4468 9045 4471
rect 8996 4440 9045 4468
rect 8996 4428 9002 4440
rect 9033 4437 9045 4440
rect 9079 4437 9091 4471
rect 9033 4431 9091 4437
rect 10502 4428 10508 4480
rect 10560 4468 10566 4480
rect 10597 4471 10655 4477
rect 10597 4468 10609 4471
rect 10560 4440 10609 4468
rect 10560 4428 10566 4440
rect 10597 4437 10609 4440
rect 10643 4437 10655 4471
rect 10597 4431 10655 4437
rect 13262 4428 13268 4480
rect 13320 4468 13326 4480
rect 13725 4471 13783 4477
rect 13725 4468 13737 4471
rect 13320 4440 13737 4468
rect 13320 4428 13326 4440
rect 13725 4437 13737 4440
rect 13771 4437 13783 4471
rect 13725 4431 13783 4437
rect 552 4378 15364 4400
rect 552 4326 2249 4378
rect 2301 4326 2313 4378
rect 2365 4326 2377 4378
rect 2429 4326 2441 4378
rect 2493 4326 2505 4378
rect 2557 4326 5951 4378
rect 6003 4326 6015 4378
rect 6067 4326 6079 4378
rect 6131 4326 6143 4378
rect 6195 4326 6207 4378
rect 6259 4326 9653 4378
rect 9705 4326 9717 4378
rect 9769 4326 9781 4378
rect 9833 4326 9845 4378
rect 9897 4326 9909 4378
rect 9961 4326 13355 4378
rect 13407 4326 13419 4378
rect 13471 4326 13483 4378
rect 13535 4326 13547 4378
rect 13599 4326 13611 4378
rect 13663 4326 15364 4378
rect 552 4304 15364 4326
rect 8202 4224 8208 4276
rect 8260 4264 8266 4276
rect 8260 4236 10456 4264
rect 8260 4224 8266 4236
rect 6362 4088 6368 4140
rect 6420 4128 6426 4140
rect 6457 4131 6515 4137
rect 6457 4128 6469 4131
rect 6420 4100 6469 4128
rect 6420 4088 6426 4100
rect 6457 4097 6469 4100
rect 6503 4128 6515 4131
rect 8573 4131 8631 4137
rect 8573 4128 8585 4131
rect 6503 4100 8585 4128
rect 6503 4097 6515 4100
rect 6457 4091 6515 4097
rect 8573 4097 8585 4100
rect 8619 4128 8631 4131
rect 8754 4128 8760 4140
rect 8619 4100 8760 4128
rect 8619 4097 8631 4100
rect 8573 4091 8631 4097
rect 8754 4088 8760 4100
rect 8812 4088 8818 4140
rect 8938 4088 8944 4140
rect 8996 4088 9002 4140
rect 10428 4128 10456 4236
rect 13078 4224 13084 4276
rect 13136 4224 13142 4276
rect 13357 4267 13415 4273
rect 13357 4233 13369 4267
rect 13403 4264 13415 4267
rect 13403 4236 13860 4264
rect 13403 4233 13415 4236
rect 13357 4227 13415 4233
rect 10502 4156 10508 4208
rect 10560 4196 10566 4208
rect 10873 4199 10931 4205
rect 10873 4196 10885 4199
rect 10560 4168 10885 4196
rect 10560 4156 10566 4168
rect 10873 4165 10885 4168
rect 10919 4165 10931 4199
rect 10873 4159 10931 4165
rect 11057 4199 11115 4205
rect 11057 4165 11069 4199
rect 11103 4196 11115 4199
rect 11238 4196 11244 4208
rect 11103 4168 11244 4196
rect 11103 4165 11115 4168
rect 11057 4159 11115 4165
rect 11238 4156 11244 4168
rect 11296 4156 11302 4208
rect 11514 4196 11520 4208
rect 11495 4168 11520 4196
rect 11514 4156 11520 4168
rect 11572 4156 11578 4208
rect 13722 4156 13728 4208
rect 13780 4156 13786 4208
rect 13832 4196 13860 4236
rect 13906 4224 13912 4276
rect 13964 4264 13970 4276
rect 14185 4267 14243 4273
rect 14185 4264 14197 4267
rect 13964 4236 14197 4264
rect 13964 4224 13970 4236
rect 14185 4233 14197 4236
rect 14231 4233 14243 4267
rect 14185 4227 14243 4233
rect 13832 4168 14412 4196
rect 10597 4131 10655 4137
rect 10597 4128 10609 4131
rect 9048 4100 9996 4128
rect 10428 4100 10609 4128
rect 7742 4020 7748 4072
rect 7800 4060 7806 4072
rect 8294 4060 8300 4072
rect 7800 4032 8300 4060
rect 7800 4020 7806 4032
rect 8294 4020 8300 4032
rect 8352 4060 8358 4072
rect 9048 4060 9076 4100
rect 8352 4032 9076 4060
rect 8352 4020 8358 4032
rect 6730 3952 6736 4004
rect 6788 3952 6794 4004
rect 9968 3992 9996 4100
rect 10597 4097 10609 4100
rect 10643 4128 10655 4131
rect 11532 4128 11560 4156
rect 10643 4100 11560 4128
rect 11609 4131 11667 4137
rect 10643 4097 10655 4100
rect 10597 4091 10655 4097
rect 11609 4097 11621 4131
rect 11655 4128 11667 4131
rect 13170 4128 13176 4140
rect 11655 4100 11928 4128
rect 11655 4097 11667 4100
rect 11609 4091 11667 4097
rect 11238 4020 11244 4072
rect 11296 4060 11302 4072
rect 11900 4069 11928 4100
rect 13004 4100 13176 4128
rect 13004 4069 13032 4100
rect 13170 4088 13176 4100
rect 13228 4088 13234 4140
rect 11701 4063 11759 4069
rect 11701 4060 11713 4063
rect 11296 4032 11713 4060
rect 11296 4020 11302 4032
rect 11701 4029 11713 4032
rect 11747 4029 11759 4063
rect 11701 4023 11759 4029
rect 11885 4063 11943 4069
rect 11885 4029 11897 4063
rect 11931 4029 11943 4063
rect 11885 4023 11943 4029
rect 12989 4063 13047 4069
rect 12989 4029 13001 4063
rect 13035 4029 13047 4063
rect 12989 4023 13047 4029
rect 13081 4063 13139 4069
rect 13081 4029 13093 4063
rect 13127 4029 13139 4063
rect 13188 4060 13216 4088
rect 13541 4063 13599 4069
rect 13541 4060 13553 4063
rect 13188 4032 13553 4060
rect 13081 4023 13139 4029
rect 13541 4029 13553 4032
rect 13587 4029 13599 4063
rect 13541 4023 13599 4029
rect 13725 4063 13783 4069
rect 13725 4029 13737 4063
rect 13771 4029 13783 4063
rect 13725 4023 13783 4029
rect 10226 3992 10232 4004
rect 9968 3978 10232 3992
rect 9982 3964 10232 3978
rect 10226 3952 10232 3964
rect 10284 3952 10290 4004
rect 11149 3995 11207 4001
rect 11149 3961 11161 3995
rect 11195 3961 11207 3995
rect 11149 3955 11207 3961
rect 9674 3884 9680 3936
rect 9732 3924 9738 3936
rect 10367 3927 10425 3933
rect 10367 3924 10379 3927
rect 9732 3896 10379 3924
rect 9732 3884 9738 3896
rect 10367 3893 10379 3896
rect 10413 3924 10425 3927
rect 10502 3924 10508 3936
rect 10413 3896 10508 3924
rect 10413 3893 10425 3896
rect 10367 3887 10425 3893
rect 10502 3884 10508 3896
rect 10560 3924 10566 3936
rect 11164 3924 11192 3955
rect 12802 3952 12808 4004
rect 12860 3992 12866 4004
rect 13096 3992 13124 4023
rect 12860 3964 13308 3992
rect 12860 3952 12866 3964
rect 10560 3896 11192 3924
rect 10560 3884 10566 3896
rect 11422 3884 11428 3936
rect 11480 3924 11486 3936
rect 11793 3927 11851 3933
rect 11793 3924 11805 3927
rect 11480 3896 11805 3924
rect 11480 3884 11486 3896
rect 11793 3893 11805 3896
rect 11839 3893 11851 3927
rect 13280 3924 13308 3964
rect 13740 3924 13768 4023
rect 13906 4020 13912 4072
rect 13964 4020 13970 4072
rect 14384 4069 14412 4168
rect 14369 4063 14427 4069
rect 14369 4029 14381 4063
rect 14415 4029 14427 4063
rect 14369 4023 14427 4029
rect 14461 4063 14519 4069
rect 14461 4029 14473 4063
rect 14507 4029 14519 4063
rect 14461 4023 14519 4029
rect 13814 3952 13820 4004
rect 13872 3992 13878 4004
rect 14476 3992 14504 4023
rect 13872 3964 14504 3992
rect 13872 3952 13878 3964
rect 13280 3896 13768 3924
rect 11793 3887 11851 3893
rect 552 3834 15520 3856
rect 552 3782 4100 3834
rect 4152 3782 4164 3834
rect 4216 3782 4228 3834
rect 4280 3782 4292 3834
rect 4344 3782 4356 3834
rect 4408 3782 7802 3834
rect 7854 3782 7866 3834
rect 7918 3782 7930 3834
rect 7982 3782 7994 3834
rect 8046 3782 8058 3834
rect 8110 3782 11504 3834
rect 11556 3782 11568 3834
rect 11620 3782 11632 3834
rect 11684 3782 11696 3834
rect 11748 3782 11760 3834
rect 11812 3782 15206 3834
rect 15258 3782 15270 3834
rect 15322 3782 15334 3834
rect 15386 3782 15398 3834
rect 15450 3782 15462 3834
rect 15514 3782 15520 3834
rect 552 3760 15520 3782
rect 6730 3680 6736 3732
rect 6788 3720 6794 3732
rect 7101 3723 7159 3729
rect 7101 3720 7113 3723
rect 6788 3692 7113 3720
rect 6788 3680 6794 3692
rect 7101 3689 7113 3692
rect 7147 3689 7159 3723
rect 7101 3683 7159 3689
rect 8202 3680 8208 3732
rect 8260 3680 8266 3732
rect 9214 3680 9220 3732
rect 9272 3680 9278 3732
rect 9674 3680 9680 3732
rect 9732 3680 9738 3732
rect 12802 3680 12808 3732
rect 12860 3680 12866 3732
rect 8297 3655 8355 3661
rect 8297 3621 8309 3655
rect 8343 3652 8355 3655
rect 9585 3655 9643 3661
rect 9585 3652 9597 3655
rect 8343 3624 9597 3652
rect 8343 3621 8355 3624
rect 8297 3615 8355 3621
rect 9585 3621 9597 3624
rect 9631 3652 9643 3655
rect 9631 3624 12756 3652
rect 9631 3621 9643 3624
rect 9585 3615 9643 3621
rect 7285 3587 7343 3593
rect 7285 3553 7297 3587
rect 7331 3584 7343 3587
rect 8570 3584 8576 3596
rect 7331 3556 7880 3584
rect 7331 3553 7343 3556
rect 7285 3547 7343 3553
rect 7852 3457 7880 3556
rect 8496 3556 8576 3584
rect 8496 3525 8524 3556
rect 8570 3544 8576 3556
rect 8628 3584 8634 3596
rect 8757 3587 8815 3593
rect 8757 3584 8769 3587
rect 8628 3556 8769 3584
rect 8628 3544 8634 3556
rect 8757 3553 8769 3556
rect 8803 3584 8815 3587
rect 9030 3584 9036 3596
rect 8803 3556 9036 3584
rect 8803 3553 8815 3556
rect 8757 3547 8815 3553
rect 9030 3544 9036 3556
rect 9088 3544 9094 3596
rect 9122 3544 9128 3596
rect 9180 3584 9186 3596
rect 9306 3584 9312 3596
rect 9180 3556 9312 3584
rect 9180 3544 9186 3556
rect 9306 3544 9312 3556
rect 9364 3584 9370 3596
rect 9364 3556 9812 3584
rect 9364 3544 9370 3556
rect 9784 3525 9812 3556
rect 11330 3544 11336 3596
rect 11388 3544 11394 3596
rect 12342 3584 12348 3596
rect 11716 3556 12348 3584
rect 8481 3519 8539 3525
rect 8481 3485 8493 3519
rect 8527 3485 8539 3519
rect 8481 3479 8539 3485
rect 9769 3519 9827 3525
rect 9769 3485 9781 3519
rect 9815 3485 9827 3519
rect 9769 3479 9827 3485
rect 11422 3476 11428 3528
rect 11480 3476 11486 3528
rect 11716 3525 11744 3556
rect 12342 3544 12348 3556
rect 12400 3584 12406 3596
rect 12621 3587 12679 3593
rect 12621 3584 12633 3587
rect 12400 3556 12633 3584
rect 12400 3544 12406 3556
rect 12621 3553 12633 3556
rect 12667 3553 12679 3587
rect 12621 3547 12679 3553
rect 11701 3519 11759 3525
rect 11701 3485 11713 3519
rect 11747 3485 11759 3519
rect 11701 3479 11759 3485
rect 12434 3476 12440 3528
rect 12492 3476 12498 3528
rect 12728 3516 12756 3624
rect 13262 3612 13268 3664
rect 13320 3612 13326 3664
rect 13998 3612 14004 3664
rect 14056 3612 14062 3664
rect 12986 3544 12992 3596
rect 13044 3544 13050 3596
rect 15010 3516 15016 3528
rect 12728 3488 15016 3516
rect 15010 3476 15016 3488
rect 15068 3476 15074 3528
rect 7837 3451 7895 3457
rect 7837 3417 7849 3451
rect 7883 3417 7895 3451
rect 7837 3411 7895 3417
rect 552 3290 15364 3312
rect 552 3238 2249 3290
rect 2301 3238 2313 3290
rect 2365 3238 2377 3290
rect 2429 3238 2441 3290
rect 2493 3238 2505 3290
rect 2557 3238 5951 3290
rect 6003 3238 6015 3290
rect 6067 3238 6079 3290
rect 6131 3238 6143 3290
rect 6195 3238 6207 3290
rect 6259 3238 9653 3290
rect 9705 3238 9717 3290
rect 9769 3238 9781 3290
rect 9833 3238 9845 3290
rect 9897 3238 9909 3290
rect 9961 3238 13355 3290
rect 13407 3238 13419 3290
rect 13471 3238 13483 3290
rect 13535 3238 13547 3290
rect 13599 3238 13611 3290
rect 13663 3238 15364 3290
rect 552 3216 15364 3238
rect 6362 3000 6368 3052
rect 6420 3000 6426 3052
rect 12342 3000 12348 3052
rect 12400 3000 12406 3052
rect 9490 2932 9496 2984
rect 9548 2972 9554 2984
rect 9677 2975 9735 2981
rect 9677 2972 9689 2975
rect 9548 2944 9689 2972
rect 9548 2932 9554 2944
rect 9677 2941 9689 2944
rect 9723 2941 9735 2975
rect 9677 2935 9735 2941
rect 12253 2975 12311 2981
rect 12253 2941 12265 2975
rect 12299 2972 12311 2975
rect 12434 2972 12440 2984
rect 12299 2944 12440 2972
rect 12299 2941 12311 2944
rect 12253 2935 12311 2941
rect 12434 2932 12440 2944
rect 12492 2932 12498 2984
rect 6638 2864 6644 2916
rect 6696 2864 6702 2916
rect 7650 2864 7656 2916
rect 7708 2864 7714 2916
rect 8113 2839 8171 2845
rect 8113 2805 8125 2839
rect 8159 2836 8171 2839
rect 8202 2836 8208 2848
rect 8159 2808 8208 2836
rect 8159 2805 8171 2808
rect 8113 2799 8171 2805
rect 8202 2796 8208 2808
rect 8260 2796 8266 2848
rect 9306 2796 9312 2848
rect 9364 2836 9370 2848
rect 9493 2839 9551 2845
rect 9493 2836 9505 2839
rect 9364 2808 9505 2836
rect 9364 2796 9370 2808
rect 9493 2805 9505 2808
rect 9539 2805 9551 2839
rect 9493 2799 9551 2805
rect 12621 2839 12679 2845
rect 12621 2805 12633 2839
rect 12667 2836 12679 2839
rect 12710 2836 12716 2848
rect 12667 2808 12716 2836
rect 12667 2805 12679 2808
rect 12621 2799 12679 2805
rect 12710 2796 12716 2808
rect 12768 2796 12774 2848
rect 552 2746 15520 2768
rect 552 2694 4100 2746
rect 4152 2694 4164 2746
rect 4216 2694 4228 2746
rect 4280 2694 4292 2746
rect 4344 2694 4356 2746
rect 4408 2694 7802 2746
rect 7854 2694 7866 2746
rect 7918 2694 7930 2746
rect 7982 2694 7994 2746
rect 8046 2694 8058 2746
rect 8110 2694 11504 2746
rect 11556 2694 11568 2746
rect 11620 2694 11632 2746
rect 11684 2694 11696 2746
rect 11748 2694 11760 2746
rect 11812 2694 15206 2746
rect 15258 2694 15270 2746
rect 15322 2694 15334 2746
rect 15386 2694 15398 2746
rect 15450 2694 15462 2746
rect 15514 2694 15520 2746
rect 552 2672 15520 2694
rect 6638 2592 6644 2644
rect 6696 2632 6702 2644
rect 7193 2635 7251 2641
rect 7193 2632 7205 2635
rect 6696 2604 7205 2632
rect 6696 2592 6702 2604
rect 7193 2601 7205 2604
rect 7239 2601 7251 2635
rect 12986 2632 12992 2644
rect 7193 2595 7251 2601
rect 9048 2604 12992 2632
rect 8202 2524 8208 2576
rect 8260 2564 8266 2576
rect 8260 2536 8708 2564
rect 8260 2524 8266 2536
rect 7377 2499 7435 2505
rect 7377 2465 7389 2499
rect 7423 2496 7435 2499
rect 7423 2468 7880 2496
rect 7423 2465 7435 2468
rect 7377 2459 7435 2465
rect 7852 2369 7880 2468
rect 8294 2456 8300 2508
rect 8352 2456 8358 2508
rect 8481 2431 8539 2437
rect 8481 2397 8493 2431
rect 8527 2428 8539 2431
rect 8680 2428 8708 2536
rect 8754 2456 8760 2508
rect 8812 2496 8818 2508
rect 8941 2499 8999 2505
rect 8941 2496 8953 2499
rect 8812 2468 8953 2496
rect 8812 2456 8818 2468
rect 8941 2465 8953 2468
rect 8987 2496 8999 2499
rect 9048 2496 9076 2604
rect 12986 2592 12992 2604
rect 13044 2592 13050 2644
rect 10318 2524 10324 2576
rect 10376 2524 10382 2576
rect 13998 2524 14004 2576
rect 14056 2524 14062 2576
rect 8987 2468 9076 2496
rect 8987 2465 8999 2468
rect 8941 2459 8999 2465
rect 9306 2456 9312 2508
rect 9364 2456 9370 2508
rect 12710 2456 12716 2508
rect 12768 2456 12774 2508
rect 12986 2456 12992 2508
rect 13044 2456 13050 2508
rect 15010 2456 15016 2508
rect 15068 2456 15074 2508
rect 10870 2428 10876 2440
rect 8527 2400 8616 2428
rect 8680 2400 10876 2428
rect 8527 2397 8539 2400
rect 8481 2391 8539 2397
rect 7837 2363 7895 2369
rect 7837 2329 7849 2363
rect 7883 2329 7895 2363
rect 7837 2323 7895 2329
rect 8588 2292 8616 2400
rect 10870 2388 10876 2400
rect 10928 2388 10934 2440
rect 12526 2388 12532 2440
rect 12584 2388 12590 2440
rect 13262 2388 13268 2440
rect 13320 2388 13326 2440
rect 9122 2292 9128 2304
rect 8588 2264 9128 2292
rect 9122 2252 9128 2264
rect 9180 2252 9186 2304
rect 10134 2252 10140 2304
rect 10192 2292 10198 2304
rect 10735 2295 10793 2301
rect 10735 2292 10747 2295
rect 10192 2264 10747 2292
rect 10192 2252 10198 2264
rect 10735 2261 10747 2264
rect 10781 2292 10793 2295
rect 11422 2292 11428 2304
rect 10781 2264 11428 2292
rect 10781 2261 10793 2264
rect 10735 2255 10793 2261
rect 11422 2252 11428 2264
rect 11480 2252 11486 2304
rect 12894 2252 12900 2304
rect 12952 2252 12958 2304
rect 552 2202 15364 2224
rect 552 2150 2249 2202
rect 2301 2150 2313 2202
rect 2365 2150 2377 2202
rect 2429 2150 2441 2202
rect 2493 2150 2505 2202
rect 2557 2150 5951 2202
rect 6003 2150 6015 2202
rect 6067 2150 6079 2202
rect 6131 2150 6143 2202
rect 6195 2150 6207 2202
rect 6259 2150 9653 2202
rect 9705 2150 9717 2202
rect 9769 2150 9781 2202
rect 9833 2150 9845 2202
rect 9897 2150 9909 2202
rect 9961 2150 13355 2202
rect 13407 2150 13419 2202
rect 13471 2150 13483 2202
rect 13535 2150 13547 2202
rect 13599 2150 13611 2202
rect 13663 2150 15364 2202
rect 552 2128 15364 2150
rect 9490 2048 9496 2100
rect 9548 2088 9554 2100
rect 9677 2091 9735 2097
rect 9677 2088 9689 2091
rect 9548 2060 9689 2088
rect 9548 2048 9554 2060
rect 9677 2057 9689 2060
rect 9723 2057 9735 2091
rect 9677 2051 9735 2057
rect 11330 2048 11336 2100
rect 11388 2088 11394 2100
rect 11425 2091 11483 2097
rect 11425 2088 11437 2091
rect 11388 2060 11437 2088
rect 11388 2048 11394 2060
rect 11425 2057 11437 2060
rect 11471 2057 11483 2091
rect 11425 2051 11483 2057
rect 13262 2048 13268 2100
rect 13320 2088 13326 2100
rect 13541 2091 13599 2097
rect 13541 2088 13553 2091
rect 13320 2060 13553 2088
rect 13320 2048 13326 2060
rect 13541 2057 13553 2060
rect 13587 2057 13599 2091
rect 13541 2051 13599 2057
rect 11146 2020 11152 2032
rect 8864 1992 11152 2020
rect 8864 1964 8892 1992
rect 11146 1980 11152 1992
rect 11204 1980 11210 2032
rect 8846 1912 8852 1964
rect 8904 1912 8910 1964
rect 9033 1955 9091 1961
rect 9033 1921 9045 1955
rect 9079 1952 9091 1955
rect 9122 1952 9128 1964
rect 9079 1924 9128 1952
rect 9079 1921 9091 1924
rect 9033 1915 9091 1921
rect 9122 1912 9128 1924
rect 9180 1912 9186 1964
rect 10134 1912 10140 1964
rect 10192 1912 10198 1964
rect 10321 1955 10379 1961
rect 10321 1921 10333 1955
rect 10367 1921 10379 1955
rect 10321 1915 10379 1921
rect 11333 1955 11391 1961
rect 11333 1921 11345 1955
rect 11379 1952 11391 1955
rect 12437 1955 12495 1961
rect 11379 1924 11652 1952
rect 11379 1921 11391 1924
rect 11333 1915 11391 1921
rect 8294 1844 8300 1896
rect 8352 1884 8358 1896
rect 8757 1887 8815 1893
rect 8757 1884 8769 1887
rect 8352 1856 8769 1884
rect 8352 1844 8358 1856
rect 8757 1853 8769 1856
rect 8803 1853 8815 1887
rect 8757 1847 8815 1853
rect 10042 1776 10048 1828
rect 10100 1776 10106 1828
rect 7650 1708 7656 1760
rect 7708 1748 7714 1760
rect 8389 1751 8447 1757
rect 8389 1748 8401 1751
rect 7708 1720 8401 1748
rect 7708 1708 7714 1720
rect 8389 1717 8401 1720
rect 8435 1717 8447 1751
rect 8389 1711 8447 1717
rect 9122 1708 9128 1760
rect 9180 1748 9186 1760
rect 10134 1748 10140 1760
rect 9180 1720 10140 1748
rect 9180 1708 9186 1720
rect 10134 1708 10140 1720
rect 10192 1748 10198 1760
rect 10336 1748 10364 1915
rect 11624 1893 11652 1924
rect 12437 1921 12449 1955
rect 12483 1952 12495 1955
rect 12526 1952 12532 1964
rect 12483 1924 12532 1952
rect 12483 1921 12495 1924
rect 12437 1915 12495 1921
rect 12526 1912 12532 1924
rect 12584 1952 12590 1964
rect 12584 1924 12848 1952
rect 12584 1912 12590 1924
rect 11609 1887 11667 1893
rect 11609 1853 11621 1887
rect 11655 1853 11667 1887
rect 11609 1847 11667 1853
rect 11885 1887 11943 1893
rect 11885 1853 11897 1887
rect 11931 1884 11943 1887
rect 11977 1887 12035 1893
rect 11977 1884 11989 1887
rect 11931 1856 11989 1884
rect 11931 1853 11943 1856
rect 11885 1847 11943 1853
rect 11977 1853 11989 1856
rect 12023 1853 12035 1887
rect 11977 1847 12035 1853
rect 10870 1776 10876 1828
rect 10928 1776 10934 1828
rect 11992 1816 12020 1847
rect 12066 1844 12072 1896
rect 12124 1884 12130 1896
rect 12253 1887 12311 1893
rect 12253 1884 12265 1887
rect 12124 1856 12265 1884
rect 12124 1844 12130 1856
rect 12253 1853 12265 1856
rect 12299 1853 12311 1887
rect 12253 1847 12311 1853
rect 12342 1844 12348 1896
rect 12400 1884 12406 1896
rect 12713 1887 12771 1893
rect 12713 1884 12725 1887
rect 12400 1856 12725 1884
rect 12400 1844 12406 1856
rect 12713 1853 12725 1856
rect 12759 1853 12771 1887
rect 12820 1884 12848 1924
rect 12894 1912 12900 1964
rect 12952 1952 12958 1964
rect 12952 1924 13584 1952
rect 12952 1912 12958 1924
rect 13078 1884 13084 1896
rect 12820 1856 13084 1884
rect 12713 1847 12771 1853
rect 13078 1844 13084 1856
rect 13136 1844 13142 1896
rect 13556 1893 13584 1924
rect 13265 1887 13323 1893
rect 13265 1853 13277 1887
rect 13311 1853 13323 1887
rect 13265 1847 13323 1853
rect 13541 1887 13599 1893
rect 13541 1853 13553 1887
rect 13587 1853 13599 1887
rect 13541 1847 13599 1853
rect 13725 1887 13783 1893
rect 13725 1853 13737 1887
rect 13771 1884 13783 1887
rect 13906 1884 13912 1896
rect 13771 1856 13912 1884
rect 13771 1853 13783 1856
rect 13725 1847 13783 1853
rect 12618 1816 12624 1828
rect 11992 1788 12624 1816
rect 12618 1776 12624 1788
rect 12676 1776 12682 1828
rect 13280 1816 13308 1847
rect 12728 1788 13308 1816
rect 12728 1760 12756 1788
rect 10192 1720 10364 1748
rect 11793 1751 11851 1757
rect 10192 1708 10198 1720
rect 11793 1717 11805 1751
rect 11839 1748 11851 1751
rect 12069 1751 12127 1757
rect 12069 1748 12081 1751
rect 11839 1720 12081 1748
rect 11839 1717 11851 1720
rect 11793 1711 11851 1717
rect 12069 1717 12081 1720
rect 12115 1748 12127 1751
rect 12342 1748 12348 1760
rect 12115 1720 12348 1748
rect 12115 1717 12127 1720
rect 12069 1711 12127 1717
rect 12342 1708 12348 1720
rect 12400 1708 12406 1760
rect 12710 1708 12716 1760
rect 12768 1708 12774 1760
rect 12802 1708 12808 1760
rect 12860 1708 12866 1760
rect 13173 1751 13231 1757
rect 13173 1717 13185 1751
rect 13219 1748 13231 1751
rect 13740 1748 13768 1847
rect 13906 1844 13912 1856
rect 13964 1844 13970 1896
rect 13219 1720 13768 1748
rect 13219 1717 13231 1720
rect 13173 1711 13231 1717
rect 552 1658 15520 1680
rect 552 1606 4100 1658
rect 4152 1606 4164 1658
rect 4216 1606 4228 1658
rect 4280 1606 4292 1658
rect 4344 1606 4356 1658
rect 4408 1606 7802 1658
rect 7854 1606 7866 1658
rect 7918 1606 7930 1658
rect 7982 1606 7994 1658
rect 8046 1606 8058 1658
rect 8110 1606 11504 1658
rect 11556 1606 11568 1658
rect 11620 1606 11632 1658
rect 11684 1606 11696 1658
rect 11748 1606 11760 1658
rect 11812 1606 15206 1658
rect 15258 1606 15270 1658
rect 15322 1606 15334 1658
rect 15386 1606 15398 1658
rect 15450 1606 15462 1658
rect 15514 1606 15520 1658
rect 552 1584 15520 1606
rect 8619 1547 8677 1553
rect 8619 1513 8631 1547
rect 8665 1544 8677 1547
rect 8846 1544 8852 1556
rect 8665 1516 8852 1544
rect 8665 1513 8677 1516
rect 8619 1507 8677 1513
rect 8846 1504 8852 1516
rect 8904 1504 8910 1556
rect 12069 1547 12127 1553
rect 9232 1516 10364 1544
rect 9232 1476 9260 1516
rect 10336 1488 10364 1516
rect 12069 1513 12081 1547
rect 12115 1544 12127 1547
rect 12342 1544 12348 1556
rect 12115 1516 12348 1544
rect 12115 1513 12127 1516
rect 12069 1507 12127 1513
rect 12342 1504 12348 1516
rect 12400 1504 12406 1556
rect 10318 1476 10324 1488
rect 8234 1448 9260 1476
rect 10258 1448 10324 1476
rect 10318 1436 10324 1448
rect 10376 1476 10382 1488
rect 10376 1448 13754 1476
rect 10376 1436 10382 1448
rect 15010 1436 15016 1488
rect 15068 1476 15074 1488
rect 15654 1476 15660 1488
rect 15068 1448 15660 1476
rect 15068 1436 15074 1448
rect 15654 1436 15660 1448
rect 15712 1436 15718 1488
rect 6825 1411 6883 1417
rect 6825 1377 6837 1411
rect 6871 1408 6883 1411
rect 6871 1380 7328 1408
rect 6871 1377 6883 1380
rect 6825 1371 6883 1377
rect 7190 1300 7196 1352
rect 7248 1300 7254 1352
rect 7300 1340 7328 1380
rect 8754 1368 8760 1420
rect 8812 1368 8818 1420
rect 10870 1368 10876 1420
rect 10928 1408 10934 1420
rect 11425 1411 11483 1417
rect 11425 1408 11437 1411
rect 10928 1380 11437 1408
rect 10928 1368 10934 1380
rect 11425 1377 11437 1380
rect 11471 1408 11483 1411
rect 12434 1408 12440 1420
rect 11471 1380 12440 1408
rect 11471 1377 11483 1380
rect 11425 1371 11483 1377
rect 12434 1368 12440 1380
rect 12492 1368 12498 1420
rect 12986 1368 12992 1420
rect 13044 1368 13050 1420
rect 8772 1340 8800 1368
rect 7300 1312 8800 1340
rect 9030 1300 9036 1352
rect 9088 1300 9094 1352
rect 11146 1300 11152 1352
rect 11204 1300 11210 1352
rect 12158 1300 12164 1352
rect 12216 1300 12222 1352
rect 13262 1300 13268 1352
rect 13320 1300 13326 1352
rect 10502 1164 10508 1216
rect 10560 1164 10566 1216
rect 12710 1164 12716 1216
rect 12768 1204 12774 1216
rect 12805 1207 12863 1213
rect 12805 1204 12817 1207
rect 12768 1176 12817 1204
rect 12768 1164 12774 1176
rect 12805 1173 12817 1176
rect 12851 1173 12863 1207
rect 12805 1167 12863 1173
rect 552 1114 15364 1136
rect 552 1062 2249 1114
rect 2301 1062 2313 1114
rect 2365 1062 2377 1114
rect 2429 1062 2441 1114
rect 2493 1062 2505 1114
rect 2557 1062 5951 1114
rect 6003 1062 6015 1114
rect 6067 1062 6079 1114
rect 6131 1062 6143 1114
rect 6195 1062 6207 1114
rect 6259 1062 9653 1114
rect 9705 1062 9717 1114
rect 9769 1062 9781 1114
rect 9833 1062 9845 1114
rect 9897 1062 9909 1114
rect 9961 1062 13355 1114
rect 13407 1062 13419 1114
rect 13471 1062 13483 1114
rect 13535 1062 13547 1114
rect 13599 1062 13611 1114
rect 13663 1062 15364 1114
rect 552 1040 15364 1062
rect 7190 960 7196 1012
rect 7248 1000 7254 1012
rect 7377 1003 7435 1009
rect 7377 1000 7389 1003
rect 7248 972 7389 1000
rect 7248 960 7254 972
rect 7377 969 7389 972
rect 7423 969 7435 1003
rect 7377 963 7435 969
rect 8570 960 8576 1012
rect 8628 960 8634 1012
rect 9030 960 9036 1012
rect 9088 1000 9094 1012
rect 9125 1003 9183 1009
rect 9125 1000 9137 1003
rect 9088 972 9137 1000
rect 9088 960 9094 972
rect 9125 969 9137 972
rect 9171 969 9183 1003
rect 9125 963 9183 969
rect 11977 1003 12035 1009
rect 11977 969 11989 1003
rect 12023 1000 12035 1003
rect 12066 1000 12072 1012
rect 12023 972 12072 1000
rect 12023 969 12035 972
rect 11977 963 12035 969
rect 12066 960 12072 972
rect 12124 960 12130 1012
rect 12437 1003 12495 1009
rect 12437 969 12449 1003
rect 12483 969 12495 1003
rect 12437 963 12495 969
rect 9585 935 9643 941
rect 9585 901 9597 935
rect 9631 901 9643 935
rect 9585 895 9643 901
rect 11885 935 11943 941
rect 11885 901 11897 935
rect 11931 932 11943 935
rect 12342 932 12348 944
rect 11931 904 12348 932
rect 11931 901 11943 904
rect 11885 895 11943 901
rect 7561 799 7619 805
rect 7561 765 7573 799
rect 7607 796 7619 799
rect 7650 796 7656 808
rect 7607 768 7656 796
rect 7607 765 7619 768
rect 7561 759 7619 765
rect 7650 756 7656 768
rect 7708 756 7714 808
rect 8386 756 8392 808
rect 8444 756 8450 808
rect 9309 799 9367 805
rect 9309 765 9321 799
rect 9355 796 9367 799
rect 9600 796 9628 895
rect 12342 892 12348 904
rect 12400 892 12406 944
rect 10042 824 10048 876
rect 10100 824 10106 876
rect 10134 824 10140 876
rect 10192 824 10198 876
rect 12069 867 12127 873
rect 12069 864 12081 867
rect 10520 836 12081 864
rect 10520 808 10548 836
rect 12069 833 12081 836
rect 12115 833 12127 867
rect 12069 827 12127 833
rect 9355 768 9628 796
rect 9953 799 10011 805
rect 9355 765 9367 768
rect 9309 759 9367 765
rect 9953 765 9965 799
rect 9999 796 10011 799
rect 10502 796 10508 808
rect 9999 768 10508 796
rect 9999 765 10011 768
rect 9953 759 10011 765
rect 10502 756 10508 768
rect 10560 756 10566 808
rect 11422 756 11428 808
rect 11480 796 11486 808
rect 11793 799 11851 805
rect 11793 796 11805 799
rect 11480 768 11805 796
rect 11480 756 11486 768
rect 11793 765 11805 768
rect 11839 765 11851 799
rect 12084 796 12112 827
rect 12158 796 12164 808
rect 12084 768 12164 796
rect 11793 759 11851 765
rect 11808 728 11836 759
rect 12158 756 12164 768
rect 12216 756 12222 808
rect 12452 728 12480 963
rect 12618 960 12624 1012
rect 12676 960 12682 1012
rect 12802 960 12808 1012
rect 12860 960 12866 1012
rect 13173 1003 13231 1009
rect 13173 969 13185 1003
rect 13219 1000 13231 1003
rect 13262 1000 13268 1012
rect 13219 972 13268 1000
rect 13219 969 13231 972
rect 13173 963 13231 969
rect 13262 960 13268 972
rect 13320 960 13326 1012
rect 12710 824 12716 876
rect 12768 824 12774 876
rect 12989 799 13047 805
rect 12989 765 13001 799
rect 13035 796 13047 799
rect 13078 796 13084 808
rect 13035 768 13084 796
rect 13035 765 13047 768
rect 12989 759 13047 765
rect 13078 756 13084 768
rect 13136 756 13142 808
rect 11808 700 12480 728
rect 552 570 15520 592
rect 552 518 4100 570
rect 4152 518 4164 570
rect 4216 518 4228 570
rect 4280 518 4292 570
rect 4344 518 4356 570
rect 4408 518 7802 570
rect 7854 518 7866 570
rect 7918 518 7930 570
rect 7982 518 7994 570
rect 8046 518 8058 570
rect 8110 518 11504 570
rect 11556 518 11568 570
rect 11620 518 11632 570
rect 11684 518 11696 570
rect 11748 518 11760 570
rect 11812 518 15206 570
rect 15258 518 15270 570
rect 15322 518 15334 570
rect 15386 518 15398 570
rect 15450 518 15462 570
rect 15514 518 15520 570
rect 552 496 15520 518
rect 8018 416 8024 468
rect 8076 456 8082 468
rect 8386 456 8392 468
rect 8076 428 8392 456
rect 8076 416 8082 428
rect 8386 416 8392 428
rect 8444 416 8450 468
<< via1 >>
rect 2249 15206 2301 15258
rect 2313 15206 2365 15258
rect 2377 15206 2429 15258
rect 2441 15206 2493 15258
rect 2505 15206 2557 15258
rect 5951 15206 6003 15258
rect 6015 15206 6067 15258
rect 6079 15206 6131 15258
rect 6143 15206 6195 15258
rect 6207 15206 6259 15258
rect 9653 15206 9705 15258
rect 9717 15206 9769 15258
rect 9781 15206 9833 15258
rect 9845 15206 9897 15258
rect 9909 15206 9961 15258
rect 13355 15206 13407 15258
rect 13419 15206 13471 15258
rect 13483 15206 13535 15258
rect 13547 15206 13599 15258
rect 13611 15206 13663 15258
rect 2688 15147 2740 15156
rect 2688 15113 2697 15147
rect 2697 15113 2731 15147
rect 2731 15113 2740 15147
rect 2688 15104 2740 15113
rect 8024 14943 8076 14952
rect 8024 14909 8033 14943
rect 8033 14909 8067 14943
rect 8067 14909 8076 14943
rect 8024 14900 8076 14909
rect 8208 14807 8260 14816
rect 8208 14773 8217 14807
rect 8217 14773 8251 14807
rect 8251 14773 8260 14807
rect 8208 14764 8260 14773
rect 4100 14662 4152 14714
rect 4164 14662 4216 14714
rect 4228 14662 4280 14714
rect 4292 14662 4344 14714
rect 4356 14662 4408 14714
rect 7802 14662 7854 14714
rect 7866 14662 7918 14714
rect 7930 14662 7982 14714
rect 7994 14662 8046 14714
rect 8058 14662 8110 14714
rect 11504 14662 11556 14714
rect 11568 14662 11620 14714
rect 11632 14662 11684 14714
rect 11696 14662 11748 14714
rect 11760 14662 11812 14714
rect 15206 14662 15258 14714
rect 15270 14662 15322 14714
rect 15334 14662 15386 14714
rect 15398 14662 15450 14714
rect 15462 14662 15514 14714
rect 15016 14263 15068 14272
rect 15016 14229 15025 14263
rect 15025 14229 15059 14263
rect 15059 14229 15068 14263
rect 15016 14220 15068 14229
rect 2249 14118 2301 14170
rect 2313 14118 2365 14170
rect 2377 14118 2429 14170
rect 2441 14118 2493 14170
rect 2505 14118 2557 14170
rect 5951 14118 6003 14170
rect 6015 14118 6067 14170
rect 6079 14118 6131 14170
rect 6143 14118 6195 14170
rect 6207 14118 6259 14170
rect 9653 14118 9705 14170
rect 9717 14118 9769 14170
rect 9781 14118 9833 14170
rect 9845 14118 9897 14170
rect 9909 14118 9961 14170
rect 13355 14118 13407 14170
rect 13419 14118 13471 14170
rect 13483 14118 13535 14170
rect 13547 14118 13599 14170
rect 13611 14118 13663 14170
rect 8208 13812 8260 13864
rect 8668 13744 8720 13796
rect 11888 13676 11940 13728
rect 4100 13574 4152 13626
rect 4164 13574 4216 13626
rect 4228 13574 4280 13626
rect 4292 13574 4344 13626
rect 4356 13574 4408 13626
rect 7802 13574 7854 13626
rect 7866 13574 7918 13626
rect 7930 13574 7982 13626
rect 7994 13574 8046 13626
rect 8058 13574 8110 13626
rect 11504 13574 11556 13626
rect 11568 13574 11620 13626
rect 11632 13574 11684 13626
rect 11696 13574 11748 13626
rect 11760 13574 11812 13626
rect 15206 13574 15258 13626
rect 15270 13574 15322 13626
rect 15334 13574 15386 13626
rect 15398 13574 15450 13626
rect 15462 13574 15514 13626
rect 8668 13472 8720 13524
rect 11888 13404 11940 13456
rect 7012 13336 7064 13388
rect 8576 13311 8628 13320
rect 8576 13277 8585 13311
rect 8585 13277 8619 13311
rect 8619 13277 8628 13311
rect 8576 13268 8628 13277
rect 10140 13379 10192 13388
rect 10140 13345 10149 13379
rect 10149 13345 10183 13379
rect 10183 13345 10192 13379
rect 10140 13336 10192 13345
rect 10968 13311 11020 13320
rect 10968 13277 10977 13311
rect 10977 13277 11011 13311
rect 11011 13277 11020 13311
rect 10968 13268 11020 13277
rect 11244 13268 11296 13320
rect 10048 13132 10100 13184
rect 12808 13175 12860 13184
rect 12808 13141 12817 13175
rect 12817 13141 12851 13175
rect 12851 13141 12860 13175
rect 12808 13132 12860 13141
rect 15016 13175 15068 13184
rect 15016 13141 15025 13175
rect 15025 13141 15059 13175
rect 15059 13141 15068 13175
rect 15016 13132 15068 13141
rect 2249 13030 2301 13082
rect 2313 13030 2365 13082
rect 2377 13030 2429 13082
rect 2441 13030 2493 13082
rect 2505 13030 2557 13082
rect 5951 13030 6003 13082
rect 6015 13030 6067 13082
rect 6079 13030 6131 13082
rect 6143 13030 6195 13082
rect 6207 13030 6259 13082
rect 9653 13030 9705 13082
rect 9717 13030 9769 13082
rect 9781 13030 9833 13082
rect 9845 13030 9897 13082
rect 9909 13030 9961 13082
rect 13355 13030 13407 13082
rect 13419 13030 13471 13082
rect 13483 13030 13535 13082
rect 13547 13030 13599 13082
rect 13611 13030 13663 13082
rect 8576 12928 8628 12980
rect 10140 12928 10192 12980
rect 9404 12792 9456 12844
rect 10232 12792 10284 12844
rect 11980 12835 12032 12844
rect 11980 12801 11989 12835
rect 11989 12801 12023 12835
rect 12023 12801 12032 12835
rect 11980 12792 12032 12801
rect 10048 12724 10100 12776
rect 10140 12724 10192 12776
rect 11244 12724 11296 12776
rect 12808 12724 12860 12776
rect 15016 12767 15068 12776
rect 15016 12733 15025 12767
rect 15025 12733 15059 12767
rect 15059 12733 15068 12767
rect 15016 12724 15068 12733
rect 14740 12656 14792 12708
rect 12256 12631 12308 12640
rect 12256 12597 12265 12631
rect 12265 12597 12299 12631
rect 12299 12597 12308 12631
rect 12256 12588 12308 12597
rect 4100 12486 4152 12538
rect 4164 12486 4216 12538
rect 4228 12486 4280 12538
rect 4292 12486 4344 12538
rect 4356 12486 4408 12538
rect 7802 12486 7854 12538
rect 7866 12486 7918 12538
rect 7930 12486 7982 12538
rect 7994 12486 8046 12538
rect 8058 12486 8110 12538
rect 11504 12486 11556 12538
rect 11568 12486 11620 12538
rect 11632 12486 11684 12538
rect 11696 12486 11748 12538
rect 11760 12486 11812 12538
rect 15206 12486 15258 12538
rect 15270 12486 15322 12538
rect 15334 12486 15386 12538
rect 15398 12486 15450 12538
rect 15462 12486 15514 12538
rect 8668 12316 8720 12368
rect 12256 12316 12308 12368
rect 7012 12291 7064 12300
rect 7012 12257 7021 12291
rect 7021 12257 7055 12291
rect 7055 12257 7064 12291
rect 7012 12248 7064 12257
rect 10048 12291 10100 12300
rect 10048 12257 10057 12291
rect 10057 12257 10091 12291
rect 10091 12257 10100 12291
rect 10048 12248 10100 12257
rect 7288 12223 7340 12232
rect 7288 12189 7297 12223
rect 7297 12189 7331 12223
rect 7331 12189 7340 12223
rect 7288 12180 7340 12189
rect 10140 12223 10192 12232
rect 10140 12189 10149 12223
rect 10149 12189 10183 12223
rect 10183 12189 10192 12223
rect 10140 12180 10192 12189
rect 10968 12180 11020 12232
rect 10508 12112 10560 12164
rect 8760 12087 8812 12096
rect 8760 12053 8769 12087
rect 8769 12053 8803 12087
rect 8803 12053 8812 12087
rect 8760 12044 8812 12053
rect 13728 12180 13780 12232
rect 14740 12223 14792 12232
rect 14740 12189 14749 12223
rect 14749 12189 14783 12223
rect 14783 12189 14792 12223
rect 14740 12180 14792 12189
rect 12992 12044 13044 12096
rect 2249 11942 2301 11994
rect 2313 11942 2365 11994
rect 2377 11942 2429 11994
rect 2441 11942 2493 11994
rect 2505 11942 2557 11994
rect 5951 11942 6003 11994
rect 6015 11942 6067 11994
rect 6079 11942 6131 11994
rect 6143 11942 6195 11994
rect 6207 11942 6259 11994
rect 9653 11942 9705 11994
rect 9717 11942 9769 11994
rect 9781 11942 9833 11994
rect 9845 11942 9897 11994
rect 9909 11942 9961 11994
rect 13355 11942 13407 11994
rect 13419 11942 13471 11994
rect 13483 11942 13535 11994
rect 13547 11942 13599 11994
rect 13611 11942 13663 11994
rect 7288 11840 7340 11892
rect 11980 11840 12032 11892
rect 8944 11704 8996 11756
rect 10232 11704 10284 11756
rect 10508 11747 10560 11756
rect 10508 11713 10517 11747
rect 10517 11713 10551 11747
rect 10551 11713 10560 11747
rect 10508 11704 10560 11713
rect 15660 11772 15712 11824
rect 8760 11679 8812 11688
rect 8760 11645 8769 11679
rect 8769 11645 8803 11679
rect 8803 11645 8812 11679
rect 8760 11636 8812 11645
rect 11152 11636 11204 11688
rect 10140 11568 10192 11620
rect 12808 11679 12860 11688
rect 12808 11645 12817 11679
rect 12817 11645 12851 11679
rect 12851 11645 12860 11679
rect 12808 11636 12860 11645
rect 8852 11543 8904 11552
rect 8852 11509 8861 11543
rect 8861 11509 8895 11543
rect 8895 11509 8904 11543
rect 8852 11500 8904 11509
rect 12624 11500 12676 11552
rect 4100 11398 4152 11450
rect 4164 11398 4216 11450
rect 4228 11398 4280 11450
rect 4292 11398 4344 11450
rect 4356 11398 4408 11450
rect 7802 11398 7854 11450
rect 7866 11398 7918 11450
rect 7930 11398 7982 11450
rect 7994 11398 8046 11450
rect 8058 11398 8110 11450
rect 11504 11398 11556 11450
rect 11568 11398 11620 11450
rect 11632 11398 11684 11450
rect 11696 11398 11748 11450
rect 11760 11398 11812 11450
rect 15206 11398 15258 11450
rect 15270 11398 15322 11450
rect 15334 11398 15386 11450
rect 15398 11398 15450 11450
rect 15462 11398 15514 11450
rect 10876 11296 10928 11348
rect 11152 11339 11204 11348
rect 11152 11305 11161 11339
rect 11161 11305 11195 11339
rect 11195 11305 11204 11339
rect 11152 11296 11204 11305
rect 8668 11228 8720 11280
rect 8852 11228 8904 11280
rect 6920 11160 6972 11212
rect 7196 11135 7248 11144
rect 7196 11101 7205 11135
rect 7205 11101 7239 11135
rect 7239 11101 7248 11135
rect 7196 11092 7248 11101
rect 9404 11135 9456 11144
rect 9404 11101 9413 11135
rect 9413 11101 9447 11135
rect 9447 11101 9456 11135
rect 9404 11092 9456 11101
rect 10140 11203 10192 11212
rect 10140 11169 10149 11203
rect 10149 11169 10183 11203
rect 10183 11169 10192 11203
rect 10140 11160 10192 11169
rect 11152 11160 11204 11212
rect 11060 11092 11112 11144
rect 13728 11228 13780 11280
rect 12072 11160 12124 11212
rect 12808 11160 12860 11212
rect 12624 11135 12676 11144
rect 12624 11101 12633 11135
rect 12633 11101 12667 11135
rect 12667 11101 12676 11135
rect 12624 11092 12676 11101
rect 12992 11135 13044 11144
rect 12992 11101 13001 11135
rect 13001 11101 13035 11135
rect 13035 11101 13044 11135
rect 12992 11092 13044 11101
rect 14924 11092 14976 11144
rect 8760 10999 8812 11008
rect 8760 10965 8769 10999
rect 8769 10965 8803 10999
rect 8803 10965 8812 10999
rect 8760 10956 8812 10965
rect 8852 10956 8904 11008
rect 10140 10956 10192 11008
rect 2249 10854 2301 10906
rect 2313 10854 2365 10906
rect 2377 10854 2429 10906
rect 2441 10854 2493 10906
rect 2505 10854 2557 10906
rect 5951 10854 6003 10906
rect 6015 10854 6067 10906
rect 6079 10854 6131 10906
rect 6143 10854 6195 10906
rect 6207 10854 6259 10906
rect 9653 10854 9705 10906
rect 9717 10854 9769 10906
rect 9781 10854 9833 10906
rect 9845 10854 9897 10906
rect 9909 10854 9961 10906
rect 13355 10854 13407 10906
rect 13419 10854 13471 10906
rect 13483 10854 13535 10906
rect 13547 10854 13599 10906
rect 13611 10854 13663 10906
rect 7196 10752 7248 10804
rect 11152 10616 11204 10668
rect 15016 10659 15068 10668
rect 15016 10625 15025 10659
rect 15025 10625 15059 10659
rect 15059 10625 15068 10659
rect 15016 10616 15068 10625
rect 8760 10548 8812 10600
rect 10876 10591 10928 10600
rect 10876 10557 10885 10591
rect 10885 10557 10919 10591
rect 10919 10557 10928 10591
rect 10876 10548 10928 10557
rect 11060 10591 11112 10600
rect 11060 10557 11069 10591
rect 11069 10557 11103 10591
rect 11103 10557 11112 10591
rect 11060 10548 11112 10557
rect 11980 10548 12032 10600
rect 12440 10591 12492 10600
rect 12440 10557 12449 10591
rect 12449 10557 12483 10591
rect 12483 10557 12492 10591
rect 12440 10548 12492 10557
rect 11336 10412 11388 10464
rect 12348 10455 12400 10464
rect 12348 10421 12357 10455
rect 12357 10421 12391 10455
rect 12391 10421 12400 10455
rect 12348 10412 12400 10421
rect 4100 10310 4152 10362
rect 4164 10310 4216 10362
rect 4228 10310 4280 10362
rect 4292 10310 4344 10362
rect 4356 10310 4408 10362
rect 7802 10310 7854 10362
rect 7866 10310 7918 10362
rect 7930 10310 7982 10362
rect 7994 10310 8046 10362
rect 8058 10310 8110 10362
rect 11504 10310 11556 10362
rect 11568 10310 11620 10362
rect 11632 10310 11684 10362
rect 11696 10310 11748 10362
rect 11760 10310 11812 10362
rect 15206 10310 15258 10362
rect 15270 10310 15322 10362
rect 15334 10310 15386 10362
rect 15398 10310 15450 10362
rect 15462 10310 15514 10362
rect 12072 10251 12124 10260
rect 12072 10217 12081 10251
rect 12081 10217 12115 10251
rect 12115 10217 12124 10251
rect 12072 10208 12124 10217
rect 12256 10251 12308 10260
rect 12256 10217 12265 10251
rect 12265 10217 12299 10251
rect 12299 10217 12308 10251
rect 12256 10208 12308 10217
rect 8668 10140 8720 10192
rect 11336 10115 11388 10124
rect 11336 10081 11345 10115
rect 11345 10081 11379 10115
rect 11379 10081 11388 10115
rect 11336 10072 11388 10081
rect 11428 10072 11480 10124
rect 11980 10115 12032 10124
rect 11980 10081 11989 10115
rect 11989 10081 12023 10115
rect 12023 10081 12032 10115
rect 11980 10072 12032 10081
rect 12348 10072 12400 10124
rect 6920 10047 6972 10056
rect 6920 10013 6929 10047
rect 6929 10013 6963 10047
rect 6963 10013 6972 10047
rect 6920 10004 6972 10013
rect 7196 10047 7248 10056
rect 7196 10013 7205 10047
rect 7205 10013 7239 10047
rect 7239 10013 7248 10047
rect 7196 10004 7248 10013
rect 12900 10047 12952 10056
rect 12900 10013 12909 10047
rect 12909 10013 12943 10047
rect 12943 10013 12952 10047
rect 12900 10004 12952 10013
rect 12440 9936 12492 9988
rect 8760 9868 8812 9920
rect 12808 9868 12860 9920
rect 13176 9868 13228 9920
rect 15016 9911 15068 9920
rect 15016 9877 15025 9911
rect 15025 9877 15059 9911
rect 15059 9877 15068 9911
rect 15016 9868 15068 9877
rect 2249 9766 2301 9818
rect 2313 9766 2365 9818
rect 2377 9766 2429 9818
rect 2441 9766 2493 9818
rect 2505 9766 2557 9818
rect 5951 9766 6003 9818
rect 6015 9766 6067 9818
rect 6079 9766 6131 9818
rect 6143 9766 6195 9818
rect 6207 9766 6259 9818
rect 9653 9766 9705 9818
rect 9717 9766 9769 9818
rect 9781 9766 9833 9818
rect 9845 9766 9897 9818
rect 9909 9766 9961 9818
rect 13355 9766 13407 9818
rect 13419 9766 13471 9818
rect 13483 9766 13535 9818
rect 13547 9766 13599 9818
rect 13611 9766 13663 9818
rect 7196 9664 7248 9716
rect 12256 9664 12308 9716
rect 12900 9707 12952 9716
rect 12900 9673 12909 9707
rect 12909 9673 12943 9707
rect 12943 9673 12952 9707
rect 12900 9664 12952 9673
rect 8944 9571 8996 9580
rect 8944 9537 8953 9571
rect 8953 9537 8987 9571
rect 8987 9537 8996 9571
rect 8944 9528 8996 9537
rect 9036 9460 9088 9512
rect 9496 9460 9548 9512
rect 12440 9460 12492 9512
rect 12532 9503 12584 9512
rect 12532 9469 12541 9503
rect 12541 9469 12575 9503
rect 12575 9469 12584 9503
rect 12532 9460 12584 9469
rect 12808 9503 12860 9512
rect 12808 9469 12817 9503
rect 12817 9469 12851 9503
rect 12851 9469 12860 9503
rect 12808 9460 12860 9469
rect 15016 9503 15068 9512
rect 15016 9469 15025 9503
rect 15025 9469 15059 9503
rect 15059 9469 15068 9503
rect 15016 9460 15068 9469
rect 7012 9392 7064 9444
rect 8760 9367 8812 9376
rect 8760 9333 8769 9367
rect 8769 9333 8803 9367
rect 8803 9333 8812 9367
rect 8760 9324 8812 9333
rect 8852 9367 8904 9376
rect 8852 9333 8861 9367
rect 8861 9333 8895 9367
rect 8895 9333 8904 9367
rect 8852 9324 8904 9333
rect 9680 9324 9732 9376
rect 12992 9324 13044 9376
rect 4100 9222 4152 9274
rect 4164 9222 4216 9274
rect 4228 9222 4280 9274
rect 4292 9222 4344 9274
rect 4356 9222 4408 9274
rect 7802 9222 7854 9274
rect 7866 9222 7918 9274
rect 7930 9222 7982 9274
rect 7994 9222 8046 9274
rect 8058 9222 8110 9274
rect 11504 9222 11556 9274
rect 11568 9222 11620 9274
rect 11632 9222 11684 9274
rect 11696 9222 11748 9274
rect 11760 9222 11812 9274
rect 15206 9222 15258 9274
rect 15270 9222 15322 9274
rect 15334 9222 15386 9274
rect 15398 9222 15450 9274
rect 15462 9222 15514 9274
rect 8852 9120 8904 9172
rect 8668 9052 8720 9104
rect 6920 8984 6972 9036
rect 7104 8984 7156 9036
rect 8760 8984 8812 9036
rect 9680 9027 9732 9036
rect 9680 8993 9689 9027
rect 9689 8993 9723 9027
rect 9723 8993 9732 9027
rect 9680 8984 9732 8993
rect 9772 9027 9824 9036
rect 9772 8993 9781 9027
rect 9781 8993 9815 9027
rect 9815 8993 9824 9027
rect 9772 8984 9824 8993
rect 10232 9027 10284 9036
rect 10232 8993 10265 9027
rect 10265 8993 10284 9027
rect 10232 8984 10284 8993
rect 10508 9027 10560 9036
rect 10508 8993 10517 9027
rect 10517 8993 10551 9027
rect 10551 8993 10560 9027
rect 10508 8984 10560 8993
rect 11428 8984 11480 9036
rect 12164 9027 12216 9036
rect 12164 8993 12173 9027
rect 12173 8993 12207 9027
rect 12207 8993 12216 9027
rect 12164 8984 12216 8993
rect 9036 8959 9088 8968
rect 9036 8925 9045 8959
rect 9045 8925 9079 8959
rect 9079 8925 9088 8959
rect 9036 8916 9088 8925
rect 9312 8916 9364 8968
rect 9404 8916 9456 8968
rect 10048 8959 10100 8968
rect 10048 8925 10057 8959
rect 10057 8925 10091 8959
rect 10091 8925 10100 8959
rect 10048 8916 10100 8925
rect 12532 9120 12584 9172
rect 13176 9052 13228 9104
rect 13728 9052 13780 9104
rect 12348 9027 12400 9036
rect 12348 8993 12357 9027
rect 12357 8993 12391 9027
rect 12391 8993 12400 9027
rect 12348 8984 12400 8993
rect 12992 9027 13044 9036
rect 12992 8993 13001 9027
rect 13001 8993 13035 9027
rect 13035 8993 13044 9027
rect 12992 8984 13044 8993
rect 15568 8916 15620 8968
rect 8576 8823 8628 8832
rect 8576 8789 8585 8823
rect 8585 8789 8619 8823
rect 8619 8789 8628 8823
rect 8576 8780 8628 8789
rect 10692 8780 10744 8832
rect 2249 8678 2301 8730
rect 2313 8678 2365 8730
rect 2377 8678 2429 8730
rect 2441 8678 2493 8730
rect 2505 8678 2557 8730
rect 5951 8678 6003 8730
rect 6015 8678 6067 8730
rect 6079 8678 6131 8730
rect 6143 8678 6195 8730
rect 6207 8678 6259 8730
rect 9653 8678 9705 8730
rect 9717 8678 9769 8730
rect 9781 8678 9833 8730
rect 9845 8678 9897 8730
rect 9909 8678 9961 8730
rect 13355 8678 13407 8730
rect 13419 8678 13471 8730
rect 13483 8678 13535 8730
rect 13547 8678 13599 8730
rect 13611 8678 13663 8730
rect 7104 8619 7156 8628
rect 7104 8585 7113 8619
rect 7113 8585 7147 8619
rect 7147 8585 7156 8619
rect 7104 8576 7156 8585
rect 10232 8576 10284 8628
rect 10876 8576 10928 8628
rect 11152 8619 11204 8628
rect 11152 8585 11161 8619
rect 11161 8585 11195 8619
rect 11195 8585 11204 8619
rect 11152 8576 11204 8585
rect 9404 8483 9456 8492
rect 9404 8449 9413 8483
rect 9413 8449 9447 8483
rect 9447 8449 9456 8483
rect 9404 8440 9456 8449
rect 8576 8372 8628 8424
rect 9036 8372 9088 8424
rect 10232 8415 10284 8424
rect 10232 8381 10241 8415
rect 10241 8381 10275 8415
rect 10275 8381 10284 8415
rect 10232 8372 10284 8381
rect 10508 8347 10560 8356
rect 10508 8313 10517 8347
rect 10517 8313 10551 8347
rect 10551 8313 10560 8347
rect 10508 8304 10560 8313
rect 10692 8483 10744 8492
rect 10692 8449 10701 8483
rect 10701 8449 10735 8483
rect 10735 8449 10744 8483
rect 10692 8440 10744 8449
rect 10876 8483 10928 8492
rect 10876 8449 10885 8483
rect 10885 8449 10919 8483
rect 10919 8449 10928 8483
rect 10876 8440 10928 8449
rect 11244 8440 11296 8492
rect 10784 8415 10836 8424
rect 10784 8381 10793 8415
rect 10793 8381 10827 8415
rect 10827 8381 10836 8415
rect 10784 8372 10836 8381
rect 12164 8483 12216 8492
rect 12164 8449 12173 8483
rect 12173 8449 12207 8483
rect 12207 8449 12216 8483
rect 12164 8440 12216 8449
rect 12348 8372 12400 8424
rect 15660 8372 15712 8424
rect 10784 8236 10836 8288
rect 12624 8279 12676 8288
rect 12624 8245 12633 8279
rect 12633 8245 12667 8279
rect 12667 8245 12676 8279
rect 12624 8236 12676 8245
rect 4100 8134 4152 8186
rect 4164 8134 4216 8186
rect 4228 8134 4280 8186
rect 4292 8134 4344 8186
rect 4356 8134 4408 8186
rect 7802 8134 7854 8186
rect 7866 8134 7918 8186
rect 7930 8134 7982 8186
rect 7994 8134 8046 8186
rect 8058 8134 8110 8186
rect 11504 8134 11556 8186
rect 11568 8134 11620 8186
rect 11632 8134 11684 8186
rect 11696 8134 11748 8186
rect 11760 8134 11812 8186
rect 15206 8134 15258 8186
rect 15270 8134 15322 8186
rect 15334 8134 15386 8186
rect 15398 8134 15450 8186
rect 15462 8134 15514 8186
rect 8668 7964 8720 8016
rect 9220 7964 9272 8016
rect 7012 7939 7064 7948
rect 7012 7905 7021 7939
rect 7021 7905 7055 7939
rect 7055 7905 7064 7939
rect 7012 7896 7064 7905
rect 10508 8032 10560 8084
rect 10876 8032 10928 8084
rect 13176 7964 13228 8016
rect 13728 7964 13780 8016
rect 15016 8007 15068 8016
rect 15016 7973 15025 8007
rect 15025 7973 15059 8007
rect 15059 7973 15068 8007
rect 15016 7964 15068 7973
rect 7288 7871 7340 7880
rect 7288 7837 7297 7871
rect 7297 7837 7331 7871
rect 7331 7837 7340 7871
rect 7288 7828 7340 7837
rect 8944 7828 8996 7880
rect 9220 7828 9272 7880
rect 10324 7871 10376 7880
rect 10324 7837 10333 7871
rect 10333 7837 10367 7871
rect 10367 7837 10376 7871
rect 10324 7828 10376 7837
rect 12992 7939 13044 7948
rect 12992 7905 13001 7939
rect 13001 7905 13035 7939
rect 13035 7905 13044 7939
rect 12992 7896 13044 7905
rect 10048 7760 10100 7812
rect 10600 7803 10652 7812
rect 10600 7769 10609 7803
rect 10609 7769 10643 7803
rect 10643 7769 10652 7803
rect 12624 7871 12676 7880
rect 12624 7837 12633 7871
rect 12633 7837 12667 7871
rect 12667 7837 12676 7871
rect 12624 7828 12676 7837
rect 10600 7760 10652 7769
rect 8944 7735 8996 7744
rect 8944 7701 8953 7735
rect 8953 7701 8987 7735
rect 8987 7701 8996 7735
rect 8944 7692 8996 7701
rect 10324 7692 10376 7744
rect 12348 7760 12400 7812
rect 2249 7590 2301 7642
rect 2313 7590 2365 7642
rect 2377 7590 2429 7642
rect 2441 7590 2493 7642
rect 2505 7590 2557 7642
rect 5951 7590 6003 7642
rect 6015 7590 6067 7642
rect 6079 7590 6131 7642
rect 6143 7590 6195 7642
rect 6207 7590 6259 7642
rect 9653 7590 9705 7642
rect 9717 7590 9769 7642
rect 9781 7590 9833 7642
rect 9845 7590 9897 7642
rect 9909 7590 9961 7642
rect 13355 7590 13407 7642
rect 13419 7590 13471 7642
rect 13483 7590 13535 7642
rect 13547 7590 13599 7642
rect 13611 7590 13663 7642
rect 7288 7488 7340 7540
rect 12808 7488 12860 7540
rect 13176 7488 13228 7540
rect 8944 7284 8996 7336
rect 9312 7327 9364 7336
rect 9312 7293 9321 7327
rect 9321 7293 9355 7327
rect 9355 7293 9364 7327
rect 9312 7284 9364 7293
rect 13268 7420 13320 7472
rect 12624 7352 12676 7404
rect 12808 7327 12860 7336
rect 12808 7293 12817 7327
rect 12817 7293 12851 7327
rect 12851 7293 12860 7327
rect 12808 7284 12860 7293
rect 9588 7216 9640 7268
rect 12900 7259 12952 7268
rect 12900 7225 12909 7259
rect 12909 7225 12943 7259
rect 12943 7225 12952 7259
rect 12900 7216 12952 7225
rect 13268 7327 13320 7336
rect 13268 7293 13277 7327
rect 13277 7293 13311 7327
rect 13311 7293 13320 7327
rect 13268 7284 13320 7293
rect 13820 7327 13872 7336
rect 13820 7293 13829 7327
rect 13829 7293 13863 7327
rect 13863 7293 13872 7327
rect 13820 7284 13872 7293
rect 9128 7191 9180 7200
rect 9128 7157 9137 7191
rect 9137 7157 9171 7191
rect 9171 7157 9180 7191
rect 9128 7148 9180 7157
rect 13728 7148 13780 7200
rect 4100 7046 4152 7098
rect 4164 7046 4216 7098
rect 4228 7046 4280 7098
rect 4292 7046 4344 7098
rect 4356 7046 4408 7098
rect 7802 7046 7854 7098
rect 7866 7046 7918 7098
rect 7930 7046 7982 7098
rect 7994 7046 8046 7098
rect 8058 7046 8110 7098
rect 11504 7046 11556 7098
rect 11568 7046 11620 7098
rect 11632 7046 11684 7098
rect 11696 7046 11748 7098
rect 11760 7046 11812 7098
rect 15206 7046 15258 7098
rect 15270 7046 15322 7098
rect 15334 7046 15386 7098
rect 15398 7046 15450 7098
rect 15462 7046 15514 7098
rect 8116 6876 8168 6928
rect 10600 6944 10652 6996
rect 9128 6851 9180 6860
rect 9128 6817 9137 6851
rect 9137 6817 9171 6851
rect 9171 6817 9180 6851
rect 9128 6808 9180 6817
rect 10876 6808 10928 6860
rect 11980 6851 12032 6860
rect 11980 6817 11989 6851
rect 11989 6817 12023 6851
rect 12023 6817 12032 6851
rect 11980 6808 12032 6817
rect 6552 6783 6604 6792
rect 6552 6749 6561 6783
rect 6561 6749 6595 6783
rect 6595 6749 6604 6783
rect 6552 6740 6604 6749
rect 6828 6783 6880 6792
rect 6828 6749 6837 6783
rect 6837 6749 6871 6783
rect 6871 6749 6880 6783
rect 6828 6740 6880 6749
rect 8760 6783 8812 6792
rect 8760 6749 8769 6783
rect 8769 6749 8803 6783
rect 8803 6749 8812 6783
rect 8760 6740 8812 6749
rect 11244 6783 11296 6792
rect 11244 6749 11253 6783
rect 11253 6749 11287 6783
rect 11287 6749 11296 6783
rect 11244 6740 11296 6749
rect 11980 6672 12032 6724
rect 12808 6808 12860 6860
rect 8300 6647 8352 6656
rect 8300 6613 8309 6647
rect 8309 6613 8343 6647
rect 8343 6613 8352 6647
rect 8300 6604 8352 6613
rect 13268 6604 13320 6656
rect 13912 6604 13964 6656
rect 2249 6502 2301 6554
rect 2313 6502 2365 6554
rect 2377 6502 2429 6554
rect 2441 6502 2493 6554
rect 2505 6502 2557 6554
rect 5951 6502 6003 6554
rect 6015 6502 6067 6554
rect 6079 6502 6131 6554
rect 6143 6502 6195 6554
rect 6207 6502 6259 6554
rect 9653 6502 9705 6554
rect 9717 6502 9769 6554
rect 9781 6502 9833 6554
rect 9845 6502 9897 6554
rect 9909 6502 9961 6554
rect 13355 6502 13407 6554
rect 13419 6502 13471 6554
rect 13483 6502 13535 6554
rect 13547 6502 13599 6554
rect 13611 6502 13663 6554
rect 6828 6400 6880 6452
rect 8116 6400 8168 6452
rect 9312 6443 9364 6452
rect 9312 6409 9321 6443
rect 9321 6409 9355 6443
rect 9355 6409 9364 6443
rect 9312 6400 9364 6409
rect 9036 6307 9088 6316
rect 9036 6273 9045 6307
rect 9045 6273 9079 6307
rect 9079 6273 9088 6307
rect 9036 6264 9088 6273
rect 9404 6264 9456 6316
rect 9220 6196 9272 6248
rect 10600 6196 10652 6248
rect 12900 6196 12952 6248
rect 8300 6128 8352 6180
rect 9588 6128 9640 6180
rect 13728 6196 13780 6248
rect 13912 6239 13964 6248
rect 13912 6205 13921 6239
rect 13921 6205 13955 6239
rect 13955 6205 13964 6239
rect 13912 6196 13964 6205
rect 13820 6128 13872 6180
rect 8392 6060 8444 6112
rect 9128 6060 9180 6112
rect 13544 6103 13596 6112
rect 13544 6069 13553 6103
rect 13553 6069 13587 6103
rect 13587 6069 13596 6103
rect 13544 6060 13596 6069
rect 4100 5958 4152 6010
rect 4164 5958 4216 6010
rect 4228 5958 4280 6010
rect 4292 5958 4344 6010
rect 4356 5958 4408 6010
rect 7802 5958 7854 6010
rect 7866 5958 7918 6010
rect 7930 5958 7982 6010
rect 7994 5958 8046 6010
rect 8058 5958 8110 6010
rect 11504 5958 11556 6010
rect 11568 5958 11620 6010
rect 11632 5958 11684 6010
rect 11696 5958 11748 6010
rect 11760 5958 11812 6010
rect 15206 5958 15258 6010
rect 15270 5958 15322 6010
rect 15334 5958 15386 6010
rect 15398 5958 15450 6010
rect 15462 5958 15514 6010
rect 9128 5899 9180 5908
rect 9128 5865 9137 5899
rect 9137 5865 9171 5899
rect 9171 5865 9180 5899
rect 9128 5856 9180 5865
rect 15016 5856 15068 5908
rect 8208 5788 8260 5840
rect 6552 5720 6604 5772
rect 7196 5695 7248 5704
rect 7196 5661 7205 5695
rect 7205 5661 7239 5695
rect 7239 5661 7248 5695
rect 7196 5652 7248 5661
rect 8760 5652 8812 5704
rect 13544 5788 13596 5840
rect 13912 5788 13964 5840
rect 9588 5763 9640 5772
rect 9588 5729 9597 5763
rect 9597 5729 9631 5763
rect 9631 5729 9640 5763
rect 9588 5720 9640 5729
rect 9404 5695 9456 5704
rect 9404 5661 9413 5695
rect 9413 5661 9447 5695
rect 9447 5661 9456 5695
rect 9404 5652 9456 5661
rect 12992 5695 13044 5704
rect 12992 5661 13001 5695
rect 13001 5661 13035 5695
rect 13035 5661 13044 5695
rect 12992 5652 13044 5661
rect 15016 5695 15068 5704
rect 15016 5661 15025 5695
rect 15025 5661 15059 5695
rect 15059 5661 15068 5695
rect 15016 5652 15068 5661
rect 11980 5584 12032 5636
rect 8852 5516 8904 5568
rect 10048 5559 10100 5568
rect 10048 5525 10057 5559
rect 10057 5525 10091 5559
rect 10091 5525 10100 5559
rect 10048 5516 10100 5525
rect 10232 5516 10284 5568
rect 2249 5414 2301 5466
rect 2313 5414 2365 5466
rect 2377 5414 2429 5466
rect 2441 5414 2493 5466
rect 2505 5414 2557 5466
rect 5951 5414 6003 5466
rect 6015 5414 6067 5466
rect 6079 5414 6131 5466
rect 6143 5414 6195 5466
rect 6207 5414 6259 5466
rect 9653 5414 9705 5466
rect 9717 5414 9769 5466
rect 9781 5414 9833 5466
rect 9845 5414 9897 5466
rect 9909 5414 9961 5466
rect 13355 5414 13407 5466
rect 13419 5414 13471 5466
rect 13483 5414 13535 5466
rect 13547 5414 13599 5466
rect 13611 5414 13663 5466
rect 7196 5312 7248 5364
rect 11244 5312 11296 5364
rect 13728 5312 13780 5364
rect 8760 5244 8812 5296
rect 12992 5244 13044 5296
rect 8852 5108 8904 5160
rect 9496 5108 9548 5160
rect 10048 5108 10100 5160
rect 11336 5151 11388 5160
rect 11336 5117 11345 5151
rect 11345 5117 11379 5151
rect 11379 5117 11388 5151
rect 11336 5108 11388 5117
rect 11428 5108 11480 5160
rect 11060 5040 11112 5092
rect 10692 4972 10744 5024
rect 12164 5151 12216 5160
rect 12164 5117 12173 5151
rect 12173 5117 12207 5151
rect 12207 5117 12216 5151
rect 12164 5108 12216 5117
rect 12808 5151 12860 5160
rect 12808 5117 12817 5151
rect 12817 5117 12851 5151
rect 12851 5117 12860 5151
rect 12808 5108 12860 5117
rect 13728 5151 13780 5160
rect 13728 5117 13737 5151
rect 13737 5117 13771 5151
rect 13771 5117 13780 5151
rect 13728 5108 13780 5117
rect 13176 5015 13228 5024
rect 13176 4981 13185 5015
rect 13185 4981 13219 5015
rect 13219 4981 13228 5015
rect 13176 4972 13228 4981
rect 4100 4870 4152 4922
rect 4164 4870 4216 4922
rect 4228 4870 4280 4922
rect 4292 4870 4344 4922
rect 4356 4870 4408 4922
rect 7802 4870 7854 4922
rect 7866 4870 7918 4922
rect 7930 4870 7982 4922
rect 7994 4870 8046 4922
rect 8058 4870 8110 4922
rect 11504 4870 11556 4922
rect 11568 4870 11620 4922
rect 11632 4870 11684 4922
rect 11696 4870 11748 4922
rect 11760 4870 11812 4922
rect 15206 4870 15258 4922
rect 15270 4870 15322 4922
rect 15334 4870 15386 4922
rect 15398 4870 15450 4922
rect 15462 4870 15514 4922
rect 10692 4768 10744 4820
rect 11336 4768 11388 4820
rect 12808 4700 12860 4752
rect 9220 4675 9272 4684
rect 9220 4641 9229 4675
rect 9229 4641 9263 4675
rect 9263 4641 9272 4675
rect 9220 4632 9272 4641
rect 10048 4632 10100 4684
rect 10232 4675 10284 4684
rect 10232 4641 10241 4675
rect 10241 4641 10275 4675
rect 10275 4641 10284 4675
rect 10232 4632 10284 4641
rect 11244 4632 11296 4684
rect 11336 4675 11388 4684
rect 11336 4641 11345 4675
rect 11345 4641 11379 4675
rect 11379 4641 11388 4675
rect 11336 4632 11388 4641
rect 11428 4675 11480 4684
rect 11428 4641 11437 4675
rect 11437 4641 11471 4675
rect 11471 4641 11480 4675
rect 11428 4632 11480 4641
rect 11520 4632 11572 4684
rect 13728 4632 13780 4684
rect 13912 4675 13964 4684
rect 13912 4641 13921 4675
rect 13921 4641 13955 4675
rect 13955 4641 13964 4675
rect 13912 4632 13964 4641
rect 11060 4564 11112 4616
rect 12164 4496 12216 4548
rect 8944 4428 8996 4480
rect 10508 4428 10560 4480
rect 13268 4428 13320 4480
rect 2249 4326 2301 4378
rect 2313 4326 2365 4378
rect 2377 4326 2429 4378
rect 2441 4326 2493 4378
rect 2505 4326 2557 4378
rect 5951 4326 6003 4378
rect 6015 4326 6067 4378
rect 6079 4326 6131 4378
rect 6143 4326 6195 4378
rect 6207 4326 6259 4378
rect 9653 4326 9705 4378
rect 9717 4326 9769 4378
rect 9781 4326 9833 4378
rect 9845 4326 9897 4378
rect 9909 4326 9961 4378
rect 13355 4326 13407 4378
rect 13419 4326 13471 4378
rect 13483 4326 13535 4378
rect 13547 4326 13599 4378
rect 13611 4326 13663 4378
rect 8208 4267 8260 4276
rect 8208 4233 8217 4267
rect 8217 4233 8251 4267
rect 8251 4233 8260 4267
rect 8208 4224 8260 4233
rect 6368 4088 6420 4140
rect 8760 4088 8812 4140
rect 8944 4131 8996 4140
rect 8944 4097 8953 4131
rect 8953 4097 8987 4131
rect 8987 4097 8996 4131
rect 8944 4088 8996 4097
rect 13084 4267 13136 4276
rect 13084 4233 13093 4267
rect 13093 4233 13127 4267
rect 13127 4233 13136 4267
rect 13084 4224 13136 4233
rect 10508 4156 10560 4208
rect 11244 4156 11296 4208
rect 11520 4199 11572 4208
rect 11520 4165 11529 4199
rect 11529 4165 11563 4199
rect 11563 4165 11572 4199
rect 11520 4156 11572 4165
rect 13728 4199 13780 4208
rect 13728 4165 13737 4199
rect 13737 4165 13771 4199
rect 13771 4165 13780 4199
rect 13728 4156 13780 4165
rect 13912 4224 13964 4276
rect 7748 4020 7800 4072
rect 8300 4020 8352 4072
rect 6736 3995 6788 4004
rect 6736 3961 6745 3995
rect 6745 3961 6779 3995
rect 6779 3961 6788 3995
rect 6736 3952 6788 3961
rect 11244 4020 11296 4072
rect 13176 4088 13228 4140
rect 10232 3952 10284 4004
rect 9680 3884 9732 3936
rect 10508 3884 10560 3936
rect 12808 3952 12860 4004
rect 11428 3884 11480 3936
rect 13912 4063 13964 4072
rect 13912 4029 13921 4063
rect 13921 4029 13955 4063
rect 13955 4029 13964 4063
rect 13912 4020 13964 4029
rect 13820 3952 13872 4004
rect 4100 3782 4152 3834
rect 4164 3782 4216 3834
rect 4228 3782 4280 3834
rect 4292 3782 4344 3834
rect 4356 3782 4408 3834
rect 7802 3782 7854 3834
rect 7866 3782 7918 3834
rect 7930 3782 7982 3834
rect 7994 3782 8046 3834
rect 8058 3782 8110 3834
rect 11504 3782 11556 3834
rect 11568 3782 11620 3834
rect 11632 3782 11684 3834
rect 11696 3782 11748 3834
rect 11760 3782 11812 3834
rect 15206 3782 15258 3834
rect 15270 3782 15322 3834
rect 15334 3782 15386 3834
rect 15398 3782 15450 3834
rect 15462 3782 15514 3834
rect 6736 3680 6788 3732
rect 8208 3723 8260 3732
rect 8208 3689 8217 3723
rect 8217 3689 8251 3723
rect 8251 3689 8260 3723
rect 8208 3680 8260 3689
rect 9220 3723 9272 3732
rect 9220 3689 9229 3723
rect 9229 3689 9263 3723
rect 9263 3689 9272 3723
rect 9220 3680 9272 3689
rect 9680 3723 9732 3732
rect 9680 3689 9689 3723
rect 9689 3689 9723 3723
rect 9723 3689 9732 3723
rect 9680 3680 9732 3689
rect 12808 3723 12860 3732
rect 12808 3689 12817 3723
rect 12817 3689 12851 3723
rect 12851 3689 12860 3723
rect 12808 3680 12860 3689
rect 8576 3544 8628 3596
rect 9036 3544 9088 3596
rect 9128 3587 9180 3596
rect 9128 3553 9137 3587
rect 9137 3553 9171 3587
rect 9171 3553 9180 3587
rect 9128 3544 9180 3553
rect 9312 3544 9364 3596
rect 11336 3587 11388 3596
rect 11336 3553 11345 3587
rect 11345 3553 11379 3587
rect 11379 3553 11388 3587
rect 11336 3544 11388 3553
rect 11428 3519 11480 3528
rect 11428 3485 11437 3519
rect 11437 3485 11471 3519
rect 11471 3485 11480 3519
rect 11428 3476 11480 3485
rect 12348 3544 12400 3596
rect 12440 3519 12492 3528
rect 12440 3485 12449 3519
rect 12449 3485 12483 3519
rect 12483 3485 12492 3519
rect 12440 3476 12492 3485
rect 13268 3655 13320 3664
rect 13268 3621 13277 3655
rect 13277 3621 13311 3655
rect 13311 3621 13320 3655
rect 13268 3612 13320 3621
rect 14004 3612 14056 3664
rect 12992 3587 13044 3596
rect 12992 3553 13001 3587
rect 13001 3553 13035 3587
rect 13035 3553 13044 3587
rect 12992 3544 13044 3553
rect 15016 3519 15068 3528
rect 15016 3485 15025 3519
rect 15025 3485 15059 3519
rect 15059 3485 15068 3519
rect 15016 3476 15068 3485
rect 2249 3238 2301 3290
rect 2313 3238 2365 3290
rect 2377 3238 2429 3290
rect 2441 3238 2493 3290
rect 2505 3238 2557 3290
rect 5951 3238 6003 3290
rect 6015 3238 6067 3290
rect 6079 3238 6131 3290
rect 6143 3238 6195 3290
rect 6207 3238 6259 3290
rect 9653 3238 9705 3290
rect 9717 3238 9769 3290
rect 9781 3238 9833 3290
rect 9845 3238 9897 3290
rect 9909 3238 9961 3290
rect 13355 3238 13407 3290
rect 13419 3238 13471 3290
rect 13483 3238 13535 3290
rect 13547 3238 13599 3290
rect 13611 3238 13663 3290
rect 6368 3043 6420 3052
rect 6368 3009 6377 3043
rect 6377 3009 6411 3043
rect 6411 3009 6420 3043
rect 6368 3000 6420 3009
rect 12348 3043 12400 3052
rect 12348 3009 12357 3043
rect 12357 3009 12391 3043
rect 12391 3009 12400 3043
rect 12348 3000 12400 3009
rect 9496 2932 9548 2984
rect 12440 2932 12492 2984
rect 6644 2907 6696 2916
rect 6644 2873 6653 2907
rect 6653 2873 6687 2907
rect 6687 2873 6696 2907
rect 6644 2864 6696 2873
rect 7656 2864 7708 2916
rect 8208 2796 8260 2848
rect 9312 2796 9364 2848
rect 12716 2796 12768 2848
rect 4100 2694 4152 2746
rect 4164 2694 4216 2746
rect 4228 2694 4280 2746
rect 4292 2694 4344 2746
rect 4356 2694 4408 2746
rect 7802 2694 7854 2746
rect 7866 2694 7918 2746
rect 7930 2694 7982 2746
rect 7994 2694 8046 2746
rect 8058 2694 8110 2746
rect 11504 2694 11556 2746
rect 11568 2694 11620 2746
rect 11632 2694 11684 2746
rect 11696 2694 11748 2746
rect 11760 2694 11812 2746
rect 15206 2694 15258 2746
rect 15270 2694 15322 2746
rect 15334 2694 15386 2746
rect 15398 2694 15450 2746
rect 15462 2694 15514 2746
rect 6644 2592 6696 2644
rect 8208 2567 8260 2576
rect 8208 2533 8217 2567
rect 8217 2533 8251 2567
rect 8251 2533 8260 2567
rect 8208 2524 8260 2533
rect 8300 2499 8352 2508
rect 8300 2465 8309 2499
rect 8309 2465 8343 2499
rect 8343 2465 8352 2499
rect 8300 2456 8352 2465
rect 8760 2456 8812 2508
rect 12992 2592 13044 2644
rect 10324 2524 10376 2576
rect 14004 2524 14056 2576
rect 9312 2499 9364 2508
rect 9312 2465 9321 2499
rect 9321 2465 9355 2499
rect 9355 2465 9364 2499
rect 9312 2456 9364 2465
rect 12716 2499 12768 2508
rect 12716 2465 12725 2499
rect 12725 2465 12759 2499
rect 12759 2465 12768 2499
rect 12716 2456 12768 2465
rect 12992 2499 13044 2508
rect 12992 2465 13001 2499
rect 13001 2465 13035 2499
rect 13035 2465 13044 2499
rect 12992 2456 13044 2465
rect 15016 2499 15068 2508
rect 15016 2465 15025 2499
rect 15025 2465 15059 2499
rect 15059 2465 15068 2499
rect 15016 2456 15068 2465
rect 10876 2388 10928 2440
rect 12532 2431 12584 2440
rect 12532 2397 12541 2431
rect 12541 2397 12575 2431
rect 12575 2397 12584 2431
rect 12532 2388 12584 2397
rect 13268 2431 13320 2440
rect 13268 2397 13277 2431
rect 13277 2397 13311 2431
rect 13311 2397 13320 2431
rect 13268 2388 13320 2397
rect 9128 2252 9180 2304
rect 10140 2252 10192 2304
rect 11428 2252 11480 2304
rect 12900 2295 12952 2304
rect 12900 2261 12909 2295
rect 12909 2261 12943 2295
rect 12943 2261 12952 2295
rect 12900 2252 12952 2261
rect 2249 2150 2301 2202
rect 2313 2150 2365 2202
rect 2377 2150 2429 2202
rect 2441 2150 2493 2202
rect 2505 2150 2557 2202
rect 5951 2150 6003 2202
rect 6015 2150 6067 2202
rect 6079 2150 6131 2202
rect 6143 2150 6195 2202
rect 6207 2150 6259 2202
rect 9653 2150 9705 2202
rect 9717 2150 9769 2202
rect 9781 2150 9833 2202
rect 9845 2150 9897 2202
rect 9909 2150 9961 2202
rect 13355 2150 13407 2202
rect 13419 2150 13471 2202
rect 13483 2150 13535 2202
rect 13547 2150 13599 2202
rect 13611 2150 13663 2202
rect 9496 2048 9548 2100
rect 11336 2048 11388 2100
rect 13268 2048 13320 2100
rect 11152 2023 11204 2032
rect 11152 1989 11161 2023
rect 11161 1989 11195 2023
rect 11195 1989 11204 2023
rect 11152 1980 11204 1989
rect 8852 1955 8904 1964
rect 8852 1921 8861 1955
rect 8861 1921 8895 1955
rect 8895 1921 8904 1955
rect 8852 1912 8904 1921
rect 9128 1912 9180 1964
rect 10140 1955 10192 1964
rect 10140 1921 10149 1955
rect 10149 1921 10183 1955
rect 10183 1921 10192 1955
rect 10140 1912 10192 1921
rect 8300 1844 8352 1896
rect 10048 1819 10100 1828
rect 10048 1785 10057 1819
rect 10057 1785 10091 1819
rect 10091 1785 10100 1819
rect 10048 1776 10100 1785
rect 7656 1708 7708 1760
rect 9128 1708 9180 1760
rect 10140 1708 10192 1760
rect 12532 1912 12584 1964
rect 10876 1819 10928 1828
rect 10876 1785 10885 1819
rect 10885 1785 10919 1819
rect 10919 1785 10928 1819
rect 10876 1776 10928 1785
rect 12072 1844 12124 1896
rect 12348 1844 12400 1896
rect 12900 1912 12952 1964
rect 13084 1887 13136 1896
rect 13084 1853 13093 1887
rect 13093 1853 13127 1887
rect 13127 1853 13136 1887
rect 13084 1844 13136 1853
rect 12624 1776 12676 1828
rect 12348 1708 12400 1760
rect 12716 1708 12768 1760
rect 12808 1751 12860 1760
rect 12808 1717 12817 1751
rect 12817 1717 12851 1751
rect 12851 1717 12860 1751
rect 12808 1708 12860 1717
rect 13912 1844 13964 1896
rect 4100 1606 4152 1658
rect 4164 1606 4216 1658
rect 4228 1606 4280 1658
rect 4292 1606 4344 1658
rect 4356 1606 4408 1658
rect 7802 1606 7854 1658
rect 7866 1606 7918 1658
rect 7930 1606 7982 1658
rect 7994 1606 8046 1658
rect 8058 1606 8110 1658
rect 11504 1606 11556 1658
rect 11568 1606 11620 1658
rect 11632 1606 11684 1658
rect 11696 1606 11748 1658
rect 11760 1606 11812 1658
rect 15206 1606 15258 1658
rect 15270 1606 15322 1658
rect 15334 1606 15386 1658
rect 15398 1606 15450 1658
rect 15462 1606 15514 1658
rect 8852 1504 8904 1556
rect 12348 1504 12400 1556
rect 10324 1436 10376 1488
rect 15016 1479 15068 1488
rect 15016 1445 15025 1479
rect 15025 1445 15059 1479
rect 15059 1445 15068 1479
rect 15016 1436 15068 1445
rect 15660 1436 15712 1488
rect 7196 1343 7248 1352
rect 7196 1309 7205 1343
rect 7205 1309 7239 1343
rect 7239 1309 7248 1343
rect 7196 1300 7248 1309
rect 8760 1411 8812 1420
rect 8760 1377 8769 1411
rect 8769 1377 8803 1411
rect 8803 1377 8812 1411
rect 8760 1368 8812 1377
rect 10876 1368 10928 1420
rect 12440 1368 12492 1420
rect 12992 1411 13044 1420
rect 12992 1377 13001 1411
rect 13001 1377 13035 1411
rect 13035 1377 13044 1411
rect 12992 1368 13044 1377
rect 9036 1343 9088 1352
rect 9036 1309 9045 1343
rect 9045 1309 9079 1343
rect 9079 1309 9088 1343
rect 9036 1300 9088 1309
rect 11152 1343 11204 1352
rect 11152 1309 11161 1343
rect 11161 1309 11195 1343
rect 11195 1309 11204 1343
rect 11152 1300 11204 1309
rect 12164 1343 12216 1352
rect 12164 1309 12173 1343
rect 12173 1309 12207 1343
rect 12207 1309 12216 1343
rect 12164 1300 12216 1309
rect 13268 1343 13320 1352
rect 13268 1309 13277 1343
rect 13277 1309 13311 1343
rect 13311 1309 13320 1343
rect 13268 1300 13320 1309
rect 10508 1207 10560 1216
rect 10508 1173 10517 1207
rect 10517 1173 10551 1207
rect 10551 1173 10560 1207
rect 10508 1164 10560 1173
rect 12716 1164 12768 1216
rect 2249 1062 2301 1114
rect 2313 1062 2365 1114
rect 2377 1062 2429 1114
rect 2441 1062 2493 1114
rect 2505 1062 2557 1114
rect 5951 1062 6003 1114
rect 6015 1062 6067 1114
rect 6079 1062 6131 1114
rect 6143 1062 6195 1114
rect 6207 1062 6259 1114
rect 9653 1062 9705 1114
rect 9717 1062 9769 1114
rect 9781 1062 9833 1114
rect 9845 1062 9897 1114
rect 9909 1062 9961 1114
rect 13355 1062 13407 1114
rect 13419 1062 13471 1114
rect 13483 1062 13535 1114
rect 13547 1062 13599 1114
rect 13611 1062 13663 1114
rect 7196 960 7248 1012
rect 8576 1003 8628 1012
rect 8576 969 8585 1003
rect 8585 969 8619 1003
rect 8619 969 8628 1003
rect 8576 960 8628 969
rect 9036 960 9088 1012
rect 12072 960 12124 1012
rect 7656 756 7708 808
rect 8392 799 8444 808
rect 8392 765 8401 799
rect 8401 765 8435 799
rect 8435 765 8444 799
rect 8392 756 8444 765
rect 12348 892 12400 944
rect 10048 867 10100 876
rect 10048 833 10057 867
rect 10057 833 10091 867
rect 10091 833 10100 867
rect 10048 824 10100 833
rect 10140 867 10192 876
rect 10140 833 10149 867
rect 10149 833 10183 867
rect 10183 833 10192 867
rect 10140 824 10192 833
rect 10508 756 10560 808
rect 11428 756 11480 808
rect 12164 799 12216 808
rect 12164 765 12173 799
rect 12173 765 12207 799
rect 12207 765 12216 799
rect 12164 756 12216 765
rect 12624 1003 12676 1012
rect 12624 969 12633 1003
rect 12633 969 12667 1003
rect 12667 969 12676 1003
rect 12624 960 12676 969
rect 12808 1003 12860 1012
rect 12808 969 12817 1003
rect 12817 969 12851 1003
rect 12851 969 12860 1003
rect 12808 960 12860 969
rect 13268 960 13320 1012
rect 12716 867 12768 876
rect 12716 833 12725 867
rect 12725 833 12759 867
rect 12759 833 12768 867
rect 12716 824 12768 833
rect 13084 756 13136 808
rect 4100 518 4152 570
rect 4164 518 4216 570
rect 4228 518 4280 570
rect 4292 518 4344 570
rect 4356 518 4408 570
rect 7802 518 7854 570
rect 7866 518 7918 570
rect 7930 518 7982 570
rect 7994 518 8046 570
rect 8058 518 8110 570
rect 11504 518 11556 570
rect 11568 518 11620 570
rect 11632 518 11684 570
rect 11696 518 11748 570
rect 11760 518 11812 570
rect 15206 518 15258 570
rect 15270 518 15322 570
rect 15334 518 15386 570
rect 15398 518 15450 570
rect 15462 518 15514 570
rect 8024 416 8076 468
rect 8392 416 8444 468
<< metal2 >>
rect 2594 15722 2650 16000
rect 7930 15722 7986 16000
rect 2594 15694 2728 15722
rect 2594 15600 2650 15694
rect 2249 15260 2557 15269
rect 2249 15258 2255 15260
rect 2311 15258 2335 15260
rect 2391 15258 2415 15260
rect 2471 15258 2495 15260
rect 2551 15258 2557 15260
rect 2311 15206 2313 15258
rect 2493 15206 2495 15258
rect 2249 15204 2255 15206
rect 2311 15204 2335 15206
rect 2391 15204 2415 15206
rect 2471 15204 2495 15206
rect 2551 15204 2557 15206
rect 2249 15195 2557 15204
rect 2700 15162 2728 15694
rect 7930 15694 8064 15722
rect 7930 15600 7986 15694
rect 5951 15260 6259 15269
rect 5951 15258 5957 15260
rect 6013 15258 6037 15260
rect 6093 15258 6117 15260
rect 6173 15258 6197 15260
rect 6253 15258 6259 15260
rect 6013 15206 6015 15258
rect 6195 15206 6197 15258
rect 5951 15204 5957 15206
rect 6013 15204 6037 15206
rect 6093 15204 6117 15206
rect 6173 15204 6197 15206
rect 6253 15204 6259 15206
rect 5951 15195 6259 15204
rect 2688 15156 2740 15162
rect 2688 15098 2740 15104
rect 8036 14958 8064 15694
rect 13266 15600 13322 16000
rect 9653 15260 9961 15269
rect 9653 15258 9659 15260
rect 9715 15258 9739 15260
rect 9795 15258 9819 15260
rect 9875 15258 9899 15260
rect 9955 15258 9961 15260
rect 9715 15206 9717 15258
rect 9897 15206 9899 15258
rect 9653 15204 9659 15206
rect 9715 15204 9739 15206
rect 9795 15204 9819 15206
rect 9875 15204 9899 15206
rect 9955 15204 9961 15206
rect 9653 15195 9961 15204
rect 8024 14952 8076 14958
rect 8024 14894 8076 14900
rect 8208 14816 8260 14822
rect 8208 14758 8260 14764
rect 4100 14716 4408 14725
rect 4100 14714 4106 14716
rect 4162 14714 4186 14716
rect 4242 14714 4266 14716
rect 4322 14714 4346 14716
rect 4402 14714 4408 14716
rect 4162 14662 4164 14714
rect 4344 14662 4346 14714
rect 4100 14660 4106 14662
rect 4162 14660 4186 14662
rect 4242 14660 4266 14662
rect 4322 14660 4346 14662
rect 4402 14660 4408 14662
rect 4100 14651 4408 14660
rect 7802 14716 8110 14725
rect 7802 14714 7808 14716
rect 7864 14714 7888 14716
rect 7944 14714 7968 14716
rect 8024 14714 8048 14716
rect 8104 14714 8110 14716
rect 7864 14662 7866 14714
rect 8046 14662 8048 14714
rect 7802 14660 7808 14662
rect 7864 14660 7888 14662
rect 7944 14660 7968 14662
rect 8024 14660 8048 14662
rect 8104 14660 8110 14662
rect 7802 14651 8110 14660
rect 2249 14172 2557 14181
rect 2249 14170 2255 14172
rect 2311 14170 2335 14172
rect 2391 14170 2415 14172
rect 2471 14170 2495 14172
rect 2551 14170 2557 14172
rect 2311 14118 2313 14170
rect 2493 14118 2495 14170
rect 2249 14116 2255 14118
rect 2311 14116 2335 14118
rect 2391 14116 2415 14118
rect 2471 14116 2495 14118
rect 2551 14116 2557 14118
rect 2249 14107 2557 14116
rect 5951 14172 6259 14181
rect 5951 14170 5957 14172
rect 6013 14170 6037 14172
rect 6093 14170 6117 14172
rect 6173 14170 6197 14172
rect 6253 14170 6259 14172
rect 6013 14118 6015 14170
rect 6195 14118 6197 14170
rect 5951 14116 5957 14118
rect 6013 14116 6037 14118
rect 6093 14116 6117 14118
rect 6173 14116 6197 14118
rect 6253 14116 6259 14118
rect 5951 14107 6259 14116
rect 8220 13870 8248 14758
rect 11504 14716 11812 14725
rect 11504 14714 11510 14716
rect 11566 14714 11590 14716
rect 11646 14714 11670 14716
rect 11726 14714 11750 14716
rect 11806 14714 11812 14716
rect 11566 14662 11568 14714
rect 11748 14662 11750 14714
rect 11504 14660 11510 14662
rect 11566 14660 11590 14662
rect 11646 14660 11670 14662
rect 11726 14660 11750 14662
rect 11806 14660 11812 14662
rect 11504 14651 11812 14660
rect 9653 14172 9961 14181
rect 9653 14170 9659 14172
rect 9715 14170 9739 14172
rect 9795 14170 9819 14172
rect 9875 14170 9899 14172
rect 9955 14170 9961 14172
rect 9715 14118 9717 14170
rect 9897 14118 9899 14170
rect 9653 14116 9659 14118
rect 9715 14116 9739 14118
rect 9795 14116 9819 14118
rect 9875 14116 9899 14118
rect 9955 14116 9961 14118
rect 9653 14107 9961 14116
rect 8208 13864 8260 13870
rect 8208 13806 8260 13812
rect 8668 13796 8720 13802
rect 8668 13738 8720 13744
rect 4100 13628 4408 13637
rect 4100 13626 4106 13628
rect 4162 13626 4186 13628
rect 4242 13626 4266 13628
rect 4322 13626 4346 13628
rect 4402 13626 4408 13628
rect 4162 13574 4164 13626
rect 4344 13574 4346 13626
rect 4100 13572 4106 13574
rect 4162 13572 4186 13574
rect 4242 13572 4266 13574
rect 4322 13572 4346 13574
rect 4402 13572 4408 13574
rect 4100 13563 4408 13572
rect 7802 13628 8110 13637
rect 7802 13626 7808 13628
rect 7864 13626 7888 13628
rect 7944 13626 7968 13628
rect 8024 13626 8048 13628
rect 8104 13626 8110 13628
rect 7864 13574 7866 13626
rect 8046 13574 8048 13626
rect 7802 13572 7808 13574
rect 7864 13572 7888 13574
rect 7944 13572 7968 13574
rect 8024 13572 8048 13574
rect 8104 13572 8110 13574
rect 7802 13563 8110 13572
rect 8680 13530 8708 13738
rect 11888 13728 11940 13734
rect 11888 13670 11940 13676
rect 11504 13628 11812 13637
rect 11504 13626 11510 13628
rect 11566 13626 11590 13628
rect 11646 13626 11670 13628
rect 11726 13626 11750 13628
rect 11806 13626 11812 13628
rect 11566 13574 11568 13626
rect 11748 13574 11750 13626
rect 11504 13572 11510 13574
rect 11566 13572 11590 13574
rect 11646 13572 11670 13574
rect 11726 13572 11750 13574
rect 11806 13572 11812 13574
rect 11504 13563 11812 13572
rect 8668 13524 8720 13530
rect 8668 13466 8720 13472
rect 7012 13388 7064 13394
rect 7012 13330 7064 13336
rect 2249 13084 2557 13093
rect 2249 13082 2255 13084
rect 2311 13082 2335 13084
rect 2391 13082 2415 13084
rect 2471 13082 2495 13084
rect 2551 13082 2557 13084
rect 2311 13030 2313 13082
rect 2493 13030 2495 13082
rect 2249 13028 2255 13030
rect 2311 13028 2335 13030
rect 2391 13028 2415 13030
rect 2471 13028 2495 13030
rect 2551 13028 2557 13030
rect 2249 13019 2557 13028
rect 5951 13084 6259 13093
rect 5951 13082 5957 13084
rect 6013 13082 6037 13084
rect 6093 13082 6117 13084
rect 6173 13082 6197 13084
rect 6253 13082 6259 13084
rect 6013 13030 6015 13082
rect 6195 13030 6197 13082
rect 5951 13028 5957 13030
rect 6013 13028 6037 13030
rect 6093 13028 6117 13030
rect 6173 13028 6197 13030
rect 6253 13028 6259 13030
rect 5951 13019 6259 13028
rect 4100 12540 4408 12549
rect 4100 12538 4106 12540
rect 4162 12538 4186 12540
rect 4242 12538 4266 12540
rect 4322 12538 4346 12540
rect 4402 12538 4408 12540
rect 4162 12486 4164 12538
rect 4344 12486 4346 12538
rect 4100 12484 4106 12486
rect 4162 12484 4186 12486
rect 4242 12484 4266 12486
rect 4322 12484 4346 12486
rect 4402 12484 4408 12486
rect 4100 12475 4408 12484
rect 7024 12306 7052 13330
rect 8576 13320 8628 13326
rect 8576 13262 8628 13268
rect 8588 12986 8616 13262
rect 8576 12980 8628 12986
rect 8576 12922 8628 12928
rect 7802 12540 8110 12549
rect 7802 12538 7808 12540
rect 7864 12538 7888 12540
rect 7944 12538 7968 12540
rect 8024 12538 8048 12540
rect 8104 12538 8110 12540
rect 7864 12486 7866 12538
rect 8046 12486 8048 12538
rect 7802 12484 7808 12486
rect 7864 12484 7888 12486
rect 7944 12484 7968 12486
rect 8024 12484 8048 12486
rect 8104 12484 8110 12486
rect 7802 12475 8110 12484
rect 8680 12374 8708 13466
rect 11900 13462 11928 13670
rect 11888 13456 11940 13462
rect 11888 13398 11940 13404
rect 10140 13388 10192 13394
rect 10140 13330 10192 13336
rect 10048 13184 10100 13190
rect 10048 13126 10100 13132
rect 9653 13084 9961 13093
rect 9653 13082 9659 13084
rect 9715 13082 9739 13084
rect 9795 13082 9819 13084
rect 9875 13082 9899 13084
rect 9955 13082 9961 13084
rect 9715 13030 9717 13082
rect 9897 13030 9899 13082
rect 9653 13028 9659 13030
rect 9715 13028 9739 13030
rect 9795 13028 9819 13030
rect 9875 13028 9899 13030
rect 9955 13028 9961 13030
rect 9653 13019 9961 13028
rect 9404 12844 9456 12850
rect 9404 12786 9456 12792
rect 8668 12368 8720 12374
rect 8668 12310 8720 12316
rect 7012 12300 7064 12306
rect 7012 12242 7064 12248
rect 7288 12232 7340 12238
rect 7288 12174 7340 12180
rect 2249 11996 2557 12005
rect 2249 11994 2255 11996
rect 2311 11994 2335 11996
rect 2391 11994 2415 11996
rect 2471 11994 2495 11996
rect 2551 11994 2557 11996
rect 2311 11942 2313 11994
rect 2493 11942 2495 11994
rect 2249 11940 2255 11942
rect 2311 11940 2335 11942
rect 2391 11940 2415 11942
rect 2471 11940 2495 11942
rect 2551 11940 2557 11942
rect 2249 11931 2557 11940
rect 5951 11996 6259 12005
rect 5951 11994 5957 11996
rect 6013 11994 6037 11996
rect 6093 11994 6117 11996
rect 6173 11994 6197 11996
rect 6253 11994 6259 11996
rect 6013 11942 6015 11994
rect 6195 11942 6197 11994
rect 5951 11940 5957 11942
rect 6013 11940 6037 11942
rect 6093 11940 6117 11942
rect 6173 11940 6197 11942
rect 6253 11940 6259 11942
rect 5951 11931 6259 11940
rect 7300 11898 7328 12174
rect 7288 11892 7340 11898
rect 7288 11834 7340 11840
rect 4100 11452 4408 11461
rect 4100 11450 4106 11452
rect 4162 11450 4186 11452
rect 4242 11450 4266 11452
rect 4322 11450 4346 11452
rect 4402 11450 4408 11452
rect 4162 11398 4164 11450
rect 4344 11398 4346 11450
rect 4100 11396 4106 11398
rect 4162 11396 4186 11398
rect 4242 11396 4266 11398
rect 4322 11396 4346 11398
rect 4402 11396 4408 11398
rect 4100 11387 4408 11396
rect 7802 11452 8110 11461
rect 7802 11450 7808 11452
rect 7864 11450 7888 11452
rect 7944 11450 7968 11452
rect 8024 11450 8048 11452
rect 8104 11450 8110 11452
rect 7864 11398 7866 11450
rect 8046 11398 8048 11450
rect 7802 11396 7808 11398
rect 7864 11396 7888 11398
rect 7944 11396 7968 11398
rect 8024 11396 8048 11398
rect 8104 11396 8110 11398
rect 7802 11387 8110 11396
rect 8680 11286 8708 12310
rect 8760 12096 8812 12102
rect 8760 12038 8812 12044
rect 8772 11694 8800 12038
rect 8944 11756 8996 11762
rect 8944 11698 8996 11704
rect 8760 11688 8812 11694
rect 8760 11630 8812 11636
rect 8668 11280 8720 11286
rect 8668 11222 8720 11228
rect 6920 11212 6972 11218
rect 6920 11154 6972 11160
rect 2249 10908 2557 10917
rect 2249 10906 2255 10908
rect 2311 10906 2335 10908
rect 2391 10906 2415 10908
rect 2471 10906 2495 10908
rect 2551 10906 2557 10908
rect 2311 10854 2313 10906
rect 2493 10854 2495 10906
rect 2249 10852 2255 10854
rect 2311 10852 2335 10854
rect 2391 10852 2415 10854
rect 2471 10852 2495 10854
rect 2551 10852 2557 10854
rect 2249 10843 2557 10852
rect 5951 10908 6259 10917
rect 5951 10906 5957 10908
rect 6013 10906 6037 10908
rect 6093 10906 6117 10908
rect 6173 10906 6197 10908
rect 6253 10906 6259 10908
rect 6013 10854 6015 10906
rect 6195 10854 6197 10906
rect 5951 10852 5957 10854
rect 6013 10852 6037 10854
rect 6093 10852 6117 10854
rect 6173 10852 6197 10854
rect 6253 10852 6259 10854
rect 5951 10843 6259 10852
rect 4100 10364 4408 10373
rect 4100 10362 4106 10364
rect 4162 10362 4186 10364
rect 4242 10362 4266 10364
rect 4322 10362 4346 10364
rect 4402 10362 4408 10364
rect 4162 10310 4164 10362
rect 4344 10310 4346 10362
rect 4100 10308 4106 10310
rect 4162 10308 4186 10310
rect 4242 10308 4266 10310
rect 4322 10308 4346 10310
rect 4402 10308 4408 10310
rect 4100 10299 4408 10308
rect 6932 10062 6960 11154
rect 7196 11144 7248 11150
rect 7196 11086 7248 11092
rect 7208 10810 7236 11086
rect 7196 10804 7248 10810
rect 7196 10746 7248 10752
rect 7802 10364 8110 10373
rect 7802 10362 7808 10364
rect 7864 10362 7888 10364
rect 7944 10362 7968 10364
rect 8024 10362 8048 10364
rect 8104 10362 8110 10364
rect 7864 10310 7866 10362
rect 8046 10310 8048 10362
rect 7802 10308 7808 10310
rect 7864 10308 7888 10310
rect 7944 10308 7968 10310
rect 8024 10308 8048 10310
rect 8104 10308 8110 10310
rect 7802 10299 8110 10308
rect 8680 10198 8708 11222
rect 8772 11098 8800 11630
rect 8852 11552 8904 11558
rect 8852 11494 8904 11500
rect 8864 11286 8892 11494
rect 8852 11280 8904 11286
rect 8852 11222 8904 11228
rect 8772 11070 8892 11098
rect 8864 11014 8892 11070
rect 8760 11008 8812 11014
rect 8760 10950 8812 10956
rect 8852 11008 8904 11014
rect 8852 10950 8904 10956
rect 8772 10606 8800 10950
rect 8760 10600 8812 10606
rect 8760 10542 8812 10548
rect 8668 10192 8720 10198
rect 8668 10134 8720 10140
rect 6920 10056 6972 10062
rect 7196 10056 7248 10062
rect 6972 10004 7052 10010
rect 6920 9998 7052 10004
rect 7196 9998 7248 10004
rect 6932 9982 7052 9998
rect 2249 9820 2557 9829
rect 2249 9818 2255 9820
rect 2311 9818 2335 9820
rect 2391 9818 2415 9820
rect 2471 9818 2495 9820
rect 2551 9818 2557 9820
rect 2311 9766 2313 9818
rect 2493 9766 2495 9818
rect 2249 9764 2255 9766
rect 2311 9764 2335 9766
rect 2391 9764 2415 9766
rect 2471 9764 2495 9766
rect 2551 9764 2557 9766
rect 2249 9755 2557 9764
rect 5951 9820 6259 9829
rect 5951 9818 5957 9820
rect 6013 9818 6037 9820
rect 6093 9818 6117 9820
rect 6173 9818 6197 9820
rect 6253 9818 6259 9820
rect 6013 9766 6015 9818
rect 6195 9766 6197 9818
rect 5951 9764 5957 9766
rect 6013 9764 6037 9766
rect 6093 9764 6117 9766
rect 6173 9764 6197 9766
rect 6253 9764 6259 9766
rect 5951 9755 6259 9764
rect 7024 9450 7052 9982
rect 7208 9722 7236 9998
rect 7196 9716 7248 9722
rect 7196 9658 7248 9664
rect 7012 9444 7064 9450
rect 7012 9386 7064 9392
rect 4100 9276 4408 9285
rect 4100 9274 4106 9276
rect 4162 9274 4186 9276
rect 4242 9274 4266 9276
rect 4322 9274 4346 9276
rect 4402 9274 4408 9276
rect 4162 9222 4164 9274
rect 4344 9222 4346 9274
rect 4100 9220 4106 9222
rect 4162 9220 4186 9222
rect 4242 9220 4266 9222
rect 4322 9220 4346 9222
rect 4402 9220 4408 9222
rect 4100 9211 4408 9220
rect 7024 9058 7052 9386
rect 7802 9276 8110 9285
rect 7802 9274 7808 9276
rect 7864 9274 7888 9276
rect 7944 9274 7968 9276
rect 8024 9274 8048 9276
rect 8104 9274 8110 9276
rect 7864 9222 7866 9274
rect 8046 9222 8048 9274
rect 7802 9220 7808 9222
rect 7864 9220 7888 9222
rect 7944 9220 7968 9222
rect 8024 9220 8048 9222
rect 8104 9220 8110 9222
rect 7802 9211 8110 9220
rect 8680 9110 8708 10134
rect 8760 9920 8812 9926
rect 8760 9862 8812 9868
rect 8772 9382 8800 9862
rect 8956 9586 8984 11698
rect 9416 11150 9444 12786
rect 10060 12782 10088 13126
rect 10152 12986 10180 13330
rect 10968 13320 11020 13326
rect 10968 13262 11020 13268
rect 11244 13320 11296 13326
rect 11244 13262 11296 13268
rect 10140 12980 10192 12986
rect 10140 12922 10192 12928
rect 10232 12844 10284 12850
rect 10232 12786 10284 12792
rect 10048 12776 10100 12782
rect 10048 12718 10100 12724
rect 10140 12776 10192 12782
rect 10140 12718 10192 12724
rect 10060 12306 10088 12718
rect 10048 12300 10100 12306
rect 10048 12242 10100 12248
rect 10152 12238 10180 12718
rect 10140 12232 10192 12238
rect 10140 12174 10192 12180
rect 9653 11996 9961 12005
rect 9653 11994 9659 11996
rect 9715 11994 9739 11996
rect 9795 11994 9819 11996
rect 9875 11994 9899 11996
rect 9955 11994 9961 11996
rect 9715 11942 9717 11994
rect 9897 11942 9899 11994
rect 9653 11940 9659 11942
rect 9715 11940 9739 11942
rect 9795 11940 9819 11942
rect 9875 11940 9899 11942
rect 9955 11940 9961 11942
rect 9653 11931 9961 11940
rect 10244 11762 10272 12786
rect 10980 12238 11008 13262
rect 11256 12782 11284 13262
rect 11244 12776 11296 12782
rect 11244 12718 11296 12724
rect 11504 12540 11812 12549
rect 11504 12538 11510 12540
rect 11566 12538 11590 12540
rect 11646 12538 11670 12540
rect 11726 12538 11750 12540
rect 11806 12538 11812 12540
rect 11566 12486 11568 12538
rect 11748 12486 11750 12538
rect 11504 12484 11510 12486
rect 11566 12484 11590 12486
rect 11646 12484 11670 12486
rect 11726 12484 11750 12486
rect 11806 12484 11812 12486
rect 11504 12475 11812 12484
rect 10968 12232 11020 12238
rect 10968 12174 11020 12180
rect 10508 12164 10560 12170
rect 10508 12106 10560 12112
rect 10520 11762 10548 12106
rect 10232 11756 10284 11762
rect 10232 11698 10284 11704
rect 10508 11756 10560 11762
rect 10508 11698 10560 11704
rect 11152 11688 11204 11694
rect 11152 11630 11204 11636
rect 10140 11620 10192 11626
rect 10140 11562 10192 11568
rect 10152 11218 10180 11562
rect 11164 11354 11192 11630
rect 11504 11452 11812 11461
rect 11504 11450 11510 11452
rect 11566 11450 11590 11452
rect 11646 11450 11670 11452
rect 11726 11450 11750 11452
rect 11806 11450 11812 11452
rect 11566 11398 11568 11450
rect 11748 11398 11750 11450
rect 11504 11396 11510 11398
rect 11566 11396 11590 11398
rect 11646 11396 11670 11398
rect 11726 11396 11750 11398
rect 11806 11396 11812 11398
rect 11504 11387 11812 11396
rect 10876 11348 10928 11354
rect 10876 11290 10928 11296
rect 11152 11348 11204 11354
rect 11152 11290 11204 11296
rect 10140 11212 10192 11218
rect 10140 11154 10192 11160
rect 9404 11144 9456 11150
rect 9404 11086 9456 11092
rect 8944 9580 8996 9586
rect 8944 9522 8996 9528
rect 8760 9376 8812 9382
rect 8760 9318 8812 9324
rect 8852 9376 8904 9382
rect 8852 9318 8904 9324
rect 6932 9042 7052 9058
rect 8668 9104 8720 9110
rect 8668 9046 8720 9052
rect 6920 9036 7052 9042
rect 6972 9030 7052 9036
rect 6920 8978 6972 8984
rect 2249 8732 2557 8741
rect 2249 8730 2255 8732
rect 2311 8730 2335 8732
rect 2391 8730 2415 8732
rect 2471 8730 2495 8732
rect 2551 8730 2557 8732
rect 2311 8678 2313 8730
rect 2493 8678 2495 8730
rect 2249 8676 2255 8678
rect 2311 8676 2335 8678
rect 2391 8676 2415 8678
rect 2471 8676 2495 8678
rect 2551 8676 2557 8678
rect 2249 8667 2557 8676
rect 5951 8732 6259 8741
rect 5951 8730 5957 8732
rect 6013 8730 6037 8732
rect 6093 8730 6117 8732
rect 6173 8730 6197 8732
rect 6253 8730 6259 8732
rect 6013 8678 6015 8730
rect 6195 8678 6197 8730
rect 5951 8676 5957 8678
rect 6013 8676 6037 8678
rect 6093 8676 6117 8678
rect 6173 8676 6197 8678
rect 6253 8676 6259 8678
rect 5951 8667 6259 8676
rect 4100 8188 4408 8197
rect 4100 8186 4106 8188
rect 4162 8186 4186 8188
rect 4242 8186 4266 8188
rect 4322 8186 4346 8188
rect 4402 8186 4408 8188
rect 4162 8134 4164 8186
rect 4344 8134 4346 8186
rect 4100 8132 4106 8134
rect 4162 8132 4186 8134
rect 4242 8132 4266 8134
rect 4322 8132 4346 8134
rect 4402 8132 4408 8134
rect 4100 8123 4408 8132
rect 7024 7954 7052 9030
rect 7104 9036 7156 9042
rect 7104 8978 7156 8984
rect 7116 8634 7144 8978
rect 8576 8832 8628 8838
rect 8576 8774 8628 8780
rect 7104 8628 7156 8634
rect 7104 8570 7156 8576
rect 8588 8430 8616 8774
rect 8576 8424 8628 8430
rect 8576 8366 8628 8372
rect 7802 8188 8110 8197
rect 7802 8186 7808 8188
rect 7864 8186 7888 8188
rect 7944 8186 7968 8188
rect 8024 8186 8048 8188
rect 8104 8186 8110 8188
rect 7864 8134 7866 8186
rect 8046 8134 8048 8186
rect 7802 8132 7808 8134
rect 7864 8132 7888 8134
rect 7944 8132 7968 8134
rect 8024 8132 8048 8134
rect 8104 8132 8110 8134
rect 7802 8123 8110 8132
rect 8680 8022 8708 9046
rect 8772 9042 8800 9318
rect 8864 9178 8892 9318
rect 8852 9172 8904 9178
rect 8852 9114 8904 9120
rect 8760 9036 8812 9042
rect 8760 8978 8812 8984
rect 8668 8016 8720 8022
rect 8668 7958 8720 7964
rect 7012 7948 7064 7954
rect 7012 7890 7064 7896
rect 8956 7886 8984 9522
rect 9036 9512 9088 9518
rect 9036 9454 9088 9460
rect 9048 8974 9076 9454
rect 9416 9058 9444 11086
rect 10152 11014 10180 11154
rect 10140 11008 10192 11014
rect 10140 10950 10192 10956
rect 9653 10908 9961 10917
rect 9653 10906 9659 10908
rect 9715 10906 9739 10908
rect 9795 10906 9819 10908
rect 9875 10906 9899 10908
rect 9955 10906 9961 10908
rect 9715 10854 9717 10906
rect 9897 10854 9899 10906
rect 9653 10852 9659 10854
rect 9715 10852 9739 10854
rect 9795 10852 9819 10854
rect 9875 10852 9899 10854
rect 9955 10852 9961 10854
rect 9653 10843 9961 10852
rect 10888 10606 10916 11290
rect 11152 11212 11204 11218
rect 11152 11154 11204 11160
rect 11060 11144 11112 11150
rect 11060 11086 11112 11092
rect 11072 10606 11100 11086
rect 11164 10674 11192 11154
rect 11152 10668 11204 10674
rect 11152 10610 11204 10616
rect 10876 10600 10928 10606
rect 10876 10542 10928 10548
rect 11060 10600 11112 10606
rect 11060 10542 11112 10548
rect 9653 9820 9961 9829
rect 9653 9818 9659 9820
rect 9715 9818 9739 9820
rect 9795 9818 9819 9820
rect 9875 9818 9899 9820
rect 9955 9818 9961 9820
rect 9715 9766 9717 9818
rect 9897 9766 9899 9818
rect 9653 9764 9659 9766
rect 9715 9764 9739 9766
rect 9795 9764 9819 9766
rect 9875 9764 9899 9766
rect 9955 9764 9961 9766
rect 9653 9755 9961 9764
rect 9496 9512 9548 9518
rect 9496 9454 9548 9460
rect 9324 9030 9444 9058
rect 9324 8974 9352 9030
rect 9036 8968 9088 8974
rect 9036 8910 9088 8916
rect 9312 8968 9364 8974
rect 9312 8910 9364 8916
rect 9404 8968 9456 8974
rect 9404 8910 9456 8916
rect 9048 8430 9076 8910
rect 9036 8424 9088 8430
rect 9036 8366 9088 8372
rect 9220 8016 9272 8022
rect 9218 7984 9220 7993
rect 9272 7984 9274 7993
rect 9218 7919 9274 7928
rect 7288 7880 7340 7886
rect 7288 7822 7340 7828
rect 8944 7880 8996 7886
rect 9220 7880 9272 7886
rect 8996 7828 9076 7834
rect 8944 7822 9076 7828
rect 9220 7822 9272 7828
rect 2249 7644 2557 7653
rect 2249 7642 2255 7644
rect 2311 7642 2335 7644
rect 2391 7642 2415 7644
rect 2471 7642 2495 7644
rect 2551 7642 2557 7644
rect 2311 7590 2313 7642
rect 2493 7590 2495 7642
rect 2249 7588 2255 7590
rect 2311 7588 2335 7590
rect 2391 7588 2415 7590
rect 2471 7588 2495 7590
rect 2551 7588 2557 7590
rect 2249 7579 2557 7588
rect 5951 7644 6259 7653
rect 5951 7642 5957 7644
rect 6013 7642 6037 7644
rect 6093 7642 6117 7644
rect 6173 7642 6197 7644
rect 6253 7642 6259 7644
rect 6013 7590 6015 7642
rect 6195 7590 6197 7642
rect 5951 7588 5957 7590
rect 6013 7588 6037 7590
rect 6093 7588 6117 7590
rect 6173 7588 6197 7590
rect 6253 7588 6259 7590
rect 5951 7579 6259 7588
rect 7300 7546 7328 7822
rect 8956 7806 9076 7822
rect 8944 7744 8996 7750
rect 8944 7686 8996 7692
rect 7288 7540 7340 7546
rect 7288 7482 7340 7488
rect 8956 7342 8984 7686
rect 8944 7336 8996 7342
rect 8944 7278 8996 7284
rect 4100 7100 4408 7109
rect 4100 7098 4106 7100
rect 4162 7098 4186 7100
rect 4242 7098 4266 7100
rect 4322 7098 4346 7100
rect 4402 7098 4408 7100
rect 4162 7046 4164 7098
rect 4344 7046 4346 7098
rect 4100 7044 4106 7046
rect 4162 7044 4186 7046
rect 4242 7044 4266 7046
rect 4322 7044 4346 7046
rect 4402 7044 4408 7046
rect 4100 7035 4408 7044
rect 7802 7100 8110 7109
rect 7802 7098 7808 7100
rect 7864 7098 7888 7100
rect 7944 7098 7968 7100
rect 8024 7098 8048 7100
rect 8104 7098 8110 7100
rect 7864 7046 7866 7098
rect 8046 7046 8048 7098
rect 7802 7044 7808 7046
rect 7864 7044 7888 7046
rect 7944 7044 7968 7046
rect 8024 7044 8048 7046
rect 8104 7044 8110 7046
rect 7802 7035 8110 7044
rect 8116 6928 8168 6934
rect 8116 6870 8168 6876
rect 6552 6792 6604 6798
rect 6552 6734 6604 6740
rect 6828 6792 6880 6798
rect 6828 6734 6880 6740
rect 2249 6556 2557 6565
rect 2249 6554 2255 6556
rect 2311 6554 2335 6556
rect 2391 6554 2415 6556
rect 2471 6554 2495 6556
rect 2551 6554 2557 6556
rect 2311 6502 2313 6554
rect 2493 6502 2495 6554
rect 2249 6500 2255 6502
rect 2311 6500 2335 6502
rect 2391 6500 2415 6502
rect 2471 6500 2495 6502
rect 2551 6500 2557 6502
rect 2249 6491 2557 6500
rect 5951 6556 6259 6565
rect 5951 6554 5957 6556
rect 6013 6554 6037 6556
rect 6093 6554 6117 6556
rect 6173 6554 6197 6556
rect 6253 6554 6259 6556
rect 6013 6502 6015 6554
rect 6195 6502 6197 6554
rect 5951 6500 5957 6502
rect 6013 6500 6037 6502
rect 6093 6500 6117 6502
rect 6173 6500 6197 6502
rect 6253 6500 6259 6502
rect 5951 6491 6259 6500
rect 4100 6012 4408 6021
rect 4100 6010 4106 6012
rect 4162 6010 4186 6012
rect 4242 6010 4266 6012
rect 4322 6010 4346 6012
rect 4402 6010 4408 6012
rect 4162 5958 4164 6010
rect 4344 5958 4346 6010
rect 4100 5956 4106 5958
rect 4162 5956 4186 5958
rect 4242 5956 4266 5958
rect 4322 5956 4346 5958
rect 4402 5956 4408 5958
rect 4100 5947 4408 5956
rect 6564 5778 6592 6734
rect 6840 6458 6868 6734
rect 8128 6458 8156 6870
rect 8760 6792 8812 6798
rect 8760 6734 8812 6740
rect 8300 6656 8352 6662
rect 8300 6598 8352 6604
rect 6828 6452 6880 6458
rect 6828 6394 6880 6400
rect 8116 6452 8168 6458
rect 8116 6394 8168 6400
rect 8128 6202 8156 6394
rect 8128 6174 8248 6202
rect 8312 6186 8340 6598
rect 7802 6012 8110 6021
rect 7802 6010 7808 6012
rect 7864 6010 7888 6012
rect 7944 6010 7968 6012
rect 8024 6010 8048 6012
rect 8104 6010 8110 6012
rect 7864 5958 7866 6010
rect 8046 5958 8048 6010
rect 7802 5956 7808 5958
rect 7864 5956 7888 5958
rect 7944 5956 7968 5958
rect 8024 5956 8048 5958
rect 8104 5956 8110 5958
rect 7802 5947 8110 5956
rect 8220 5846 8248 6174
rect 8300 6180 8352 6186
rect 8300 6122 8352 6128
rect 8392 6112 8444 6118
rect 8392 6054 8444 6060
rect 8208 5840 8260 5846
rect 8404 5817 8432 6054
rect 8208 5782 8260 5788
rect 8390 5808 8446 5817
rect 6552 5772 6604 5778
rect 6552 5714 6604 5720
rect 7196 5704 7248 5710
rect 7196 5646 7248 5652
rect 2249 5468 2557 5477
rect 2249 5466 2255 5468
rect 2311 5466 2335 5468
rect 2391 5466 2415 5468
rect 2471 5466 2495 5468
rect 2551 5466 2557 5468
rect 2311 5414 2313 5466
rect 2493 5414 2495 5466
rect 2249 5412 2255 5414
rect 2311 5412 2335 5414
rect 2391 5412 2415 5414
rect 2471 5412 2495 5414
rect 2551 5412 2557 5414
rect 2249 5403 2557 5412
rect 5951 5468 6259 5477
rect 5951 5466 5957 5468
rect 6013 5466 6037 5468
rect 6093 5466 6117 5468
rect 6173 5466 6197 5468
rect 6253 5466 6259 5468
rect 6013 5414 6015 5466
rect 6195 5414 6197 5466
rect 5951 5412 5957 5414
rect 6013 5412 6037 5414
rect 6093 5412 6117 5414
rect 6173 5412 6197 5414
rect 6253 5412 6259 5414
rect 5951 5403 6259 5412
rect 7208 5370 7236 5646
rect 8220 5534 8248 5782
rect 8390 5743 8446 5752
rect 8772 5710 8800 6734
rect 9048 6322 9076 7806
rect 9128 7200 9180 7206
rect 9128 7142 9180 7148
rect 9140 6866 9168 7142
rect 9232 6905 9260 7822
rect 9324 7426 9352 8910
rect 9416 8498 9444 8910
rect 9404 8492 9456 8498
rect 9404 8434 9456 8440
rect 9508 7562 9536 9454
rect 9680 9376 9732 9382
rect 9680 9318 9732 9324
rect 9692 9042 9720 9318
rect 9770 9072 9826 9081
rect 9680 9036 9732 9042
rect 10506 9072 10562 9081
rect 9770 9007 9772 9016
rect 9680 8978 9732 8984
rect 9824 9007 9826 9016
rect 10232 9036 10284 9042
rect 9772 8978 9824 8984
rect 10506 9007 10508 9016
rect 10232 8978 10284 8984
rect 10560 9007 10562 9016
rect 10508 8978 10560 8984
rect 10048 8968 10100 8974
rect 10048 8910 10100 8916
rect 9653 8732 9961 8741
rect 9653 8730 9659 8732
rect 9715 8730 9739 8732
rect 9795 8730 9819 8732
rect 9875 8730 9899 8732
rect 9955 8730 9961 8732
rect 9715 8678 9717 8730
rect 9897 8678 9899 8730
rect 9653 8676 9659 8678
rect 9715 8676 9739 8678
rect 9795 8676 9819 8678
rect 9875 8676 9899 8678
rect 9955 8676 9961 8678
rect 9653 8667 9961 8676
rect 10060 7818 10088 8910
rect 10244 8786 10272 8978
rect 10692 8832 10744 8838
rect 10244 8758 10364 8786
rect 10692 8774 10744 8780
rect 10232 8628 10284 8634
rect 10232 8570 10284 8576
rect 10244 8430 10272 8570
rect 10232 8424 10284 8430
rect 10232 8366 10284 8372
rect 10336 7886 10364 8758
rect 10704 8498 10732 8774
rect 11164 8634 11192 10610
rect 11336 10464 11388 10470
rect 11336 10406 11388 10412
rect 11348 10130 11376 10406
rect 11504 10364 11812 10373
rect 11504 10362 11510 10364
rect 11566 10362 11590 10364
rect 11646 10362 11670 10364
rect 11726 10362 11750 10364
rect 11806 10362 11812 10364
rect 11566 10310 11568 10362
rect 11748 10310 11750 10362
rect 11504 10308 11510 10310
rect 11566 10308 11590 10310
rect 11646 10308 11670 10310
rect 11726 10308 11750 10310
rect 11806 10308 11812 10310
rect 11504 10299 11812 10308
rect 11336 10124 11388 10130
rect 11336 10066 11388 10072
rect 11428 10124 11480 10130
rect 11428 10066 11480 10072
rect 11440 9042 11468 10066
rect 11504 9276 11812 9285
rect 11504 9274 11510 9276
rect 11566 9274 11590 9276
rect 11646 9274 11670 9276
rect 11726 9274 11750 9276
rect 11806 9274 11812 9276
rect 11566 9222 11568 9274
rect 11748 9222 11750 9274
rect 11504 9220 11510 9222
rect 11566 9220 11590 9222
rect 11646 9220 11670 9222
rect 11726 9220 11750 9222
rect 11806 9220 11812 9222
rect 11504 9211 11812 9220
rect 11428 9036 11480 9042
rect 11428 8978 11480 8984
rect 10876 8628 10928 8634
rect 10876 8570 10928 8576
rect 11152 8628 11204 8634
rect 11152 8570 11204 8576
rect 10888 8498 10916 8570
rect 10692 8492 10744 8498
rect 10692 8434 10744 8440
rect 10876 8492 10928 8498
rect 10876 8434 10928 8440
rect 11244 8492 11296 8498
rect 11244 8434 11296 8440
rect 10784 8424 10836 8430
rect 10784 8366 10836 8372
rect 10508 8356 10560 8362
rect 10508 8298 10560 8304
rect 10520 8090 10548 8298
rect 10796 8294 10824 8366
rect 10784 8288 10836 8294
rect 10784 8230 10836 8236
rect 10796 8106 10824 8230
rect 10796 8090 10916 8106
rect 10508 8084 10560 8090
rect 10796 8084 10928 8090
rect 10796 8078 10876 8084
rect 10508 8026 10560 8032
rect 10876 8026 10928 8032
rect 10324 7880 10376 7886
rect 10324 7822 10376 7828
rect 10048 7812 10100 7818
rect 10048 7754 10100 7760
rect 10336 7750 10364 7822
rect 10600 7812 10652 7818
rect 10600 7754 10652 7760
rect 10324 7744 10376 7750
rect 10324 7686 10376 7692
rect 9653 7644 9961 7653
rect 9653 7642 9659 7644
rect 9715 7642 9739 7644
rect 9795 7642 9819 7644
rect 9875 7642 9899 7644
rect 9955 7642 9961 7644
rect 9715 7590 9717 7642
rect 9897 7590 9899 7642
rect 9653 7588 9659 7590
rect 9715 7588 9739 7590
rect 9795 7588 9819 7590
rect 9875 7588 9899 7590
rect 9955 7588 9961 7590
rect 9653 7579 9961 7588
rect 9508 7534 9628 7562
rect 9324 7398 9444 7426
rect 9312 7336 9364 7342
rect 9312 7278 9364 7284
rect 9218 6896 9274 6905
rect 9128 6860 9180 6866
rect 9218 6831 9274 6840
rect 9128 6802 9180 6808
rect 9036 6316 9088 6322
rect 9036 6258 9088 6264
rect 8760 5704 8812 5710
rect 8760 5646 8812 5652
rect 8220 5506 8340 5534
rect 7196 5364 7248 5370
rect 7196 5306 7248 5312
rect 4100 4924 4408 4933
rect 4100 4922 4106 4924
rect 4162 4922 4186 4924
rect 4242 4922 4266 4924
rect 4322 4922 4346 4924
rect 4402 4922 4408 4924
rect 4162 4870 4164 4922
rect 4344 4870 4346 4922
rect 4100 4868 4106 4870
rect 4162 4868 4186 4870
rect 4242 4868 4266 4870
rect 4322 4868 4346 4870
rect 4402 4868 4408 4870
rect 4100 4859 4408 4868
rect 7802 4924 8110 4933
rect 7802 4922 7808 4924
rect 7864 4922 7888 4924
rect 7944 4922 7968 4924
rect 8024 4922 8048 4924
rect 8104 4922 8110 4924
rect 7864 4870 7866 4922
rect 8046 4870 8048 4922
rect 7802 4868 7808 4870
rect 7864 4868 7888 4870
rect 7944 4868 7968 4870
rect 8024 4868 8048 4870
rect 8104 4868 8110 4870
rect 7802 4859 8110 4868
rect 2249 4380 2557 4389
rect 2249 4378 2255 4380
rect 2311 4378 2335 4380
rect 2391 4378 2415 4380
rect 2471 4378 2495 4380
rect 2551 4378 2557 4380
rect 2311 4326 2313 4378
rect 2493 4326 2495 4378
rect 2249 4324 2255 4326
rect 2311 4324 2335 4326
rect 2391 4324 2415 4326
rect 2471 4324 2495 4326
rect 2551 4324 2557 4326
rect 2249 4315 2557 4324
rect 5951 4380 6259 4389
rect 5951 4378 5957 4380
rect 6013 4378 6037 4380
rect 6093 4378 6117 4380
rect 6173 4378 6197 4380
rect 6253 4378 6259 4380
rect 6013 4326 6015 4378
rect 6195 4326 6197 4378
rect 5951 4324 5957 4326
rect 6013 4324 6037 4326
rect 6093 4324 6117 4326
rect 6173 4324 6197 4326
rect 6253 4324 6259 4326
rect 5951 4315 6259 4324
rect 8208 4276 8260 4282
rect 8208 4218 8260 4224
rect 6368 4140 6420 4146
rect 6368 4082 6420 4088
rect 4100 3836 4408 3845
rect 4100 3834 4106 3836
rect 4162 3834 4186 3836
rect 4242 3834 4266 3836
rect 4322 3834 4346 3836
rect 4402 3834 4408 3836
rect 4162 3782 4164 3834
rect 4344 3782 4346 3834
rect 4100 3780 4106 3782
rect 4162 3780 4186 3782
rect 4242 3780 4266 3782
rect 4322 3780 4346 3782
rect 4402 3780 4408 3782
rect 4100 3771 4408 3780
rect 2249 3292 2557 3301
rect 2249 3290 2255 3292
rect 2311 3290 2335 3292
rect 2391 3290 2415 3292
rect 2471 3290 2495 3292
rect 2551 3290 2557 3292
rect 2311 3238 2313 3290
rect 2493 3238 2495 3290
rect 2249 3236 2255 3238
rect 2311 3236 2335 3238
rect 2391 3236 2415 3238
rect 2471 3236 2495 3238
rect 2551 3236 2557 3238
rect 2249 3227 2557 3236
rect 5951 3292 6259 3301
rect 5951 3290 5957 3292
rect 6013 3290 6037 3292
rect 6093 3290 6117 3292
rect 6173 3290 6197 3292
rect 6253 3290 6259 3292
rect 6013 3238 6015 3290
rect 6195 3238 6197 3290
rect 5951 3236 5957 3238
rect 6013 3236 6037 3238
rect 6093 3236 6117 3238
rect 6173 3236 6197 3238
rect 6253 3236 6259 3238
rect 5951 3227 6259 3236
rect 6380 3058 6408 4082
rect 7748 4072 7800 4078
rect 7668 4020 7748 4026
rect 7668 4014 7800 4020
rect 6736 4004 6788 4010
rect 6736 3946 6788 3952
rect 7668 3998 7788 4014
rect 6748 3738 6776 3946
rect 6736 3732 6788 3738
rect 6736 3674 6788 3680
rect 6368 3052 6420 3058
rect 6368 2994 6420 3000
rect 7668 2922 7696 3998
rect 7802 3836 8110 3845
rect 7802 3834 7808 3836
rect 7864 3834 7888 3836
rect 7944 3834 7968 3836
rect 8024 3834 8048 3836
rect 8104 3834 8110 3836
rect 7864 3782 7866 3834
rect 8046 3782 8048 3834
rect 7802 3780 7808 3782
rect 7864 3780 7888 3782
rect 7944 3780 7968 3782
rect 8024 3780 8048 3782
rect 8104 3780 8110 3782
rect 7802 3771 8110 3780
rect 8220 3738 8248 4218
rect 8312 4078 8340 5506
rect 8772 5302 8800 5646
rect 8852 5568 8904 5574
rect 8852 5510 8904 5516
rect 8760 5296 8812 5302
rect 8760 5238 8812 5244
rect 8772 4146 8800 5238
rect 8864 5166 8892 5510
rect 8852 5160 8904 5166
rect 8852 5102 8904 5108
rect 8944 4480 8996 4486
rect 8944 4422 8996 4428
rect 8956 4146 8984 4422
rect 8760 4140 8812 4146
rect 8760 4082 8812 4088
rect 8944 4140 8996 4146
rect 8944 4082 8996 4088
rect 8300 4072 8352 4078
rect 8300 4014 8352 4020
rect 8208 3732 8260 3738
rect 8208 3674 8260 3680
rect 9048 3602 9076 6258
rect 9232 6254 9260 6831
rect 9324 6458 9352 7278
rect 9312 6452 9364 6458
rect 9312 6394 9364 6400
rect 9416 6322 9444 7398
rect 9600 7274 9628 7534
rect 9588 7268 9640 7274
rect 9588 7210 9640 7216
rect 9600 6746 9628 7210
rect 10612 7002 10640 7754
rect 10600 6996 10652 7002
rect 10600 6938 10652 6944
rect 9508 6718 9628 6746
rect 9404 6316 9456 6322
rect 9404 6258 9456 6264
rect 9220 6248 9272 6254
rect 9220 6190 9272 6196
rect 9128 6112 9180 6118
rect 9128 6054 9180 6060
rect 9140 5914 9168 6054
rect 9128 5908 9180 5914
rect 9128 5850 9180 5856
rect 9416 5710 9444 6258
rect 9404 5704 9456 5710
rect 9404 5646 9456 5652
rect 9416 5534 9444 5646
rect 9324 5506 9444 5534
rect 9220 4684 9272 4690
rect 9220 4626 9272 4632
rect 9232 3738 9260 4626
rect 9220 3732 9272 3738
rect 9220 3674 9272 3680
rect 9324 3602 9352 5506
rect 9508 5166 9536 6718
rect 9653 6556 9961 6565
rect 9653 6554 9659 6556
rect 9715 6554 9739 6556
rect 9795 6554 9819 6556
rect 9875 6554 9899 6556
rect 9955 6554 9961 6556
rect 9715 6502 9717 6554
rect 9897 6502 9899 6554
rect 9653 6500 9659 6502
rect 9715 6500 9739 6502
rect 9795 6500 9819 6502
rect 9875 6500 9899 6502
rect 9955 6500 9961 6502
rect 9653 6491 9961 6500
rect 10612 6254 10640 6938
rect 10888 6866 10916 8026
rect 10876 6860 10928 6866
rect 10876 6802 10928 6808
rect 11256 6798 11284 8434
rect 11504 8188 11812 8197
rect 11504 8186 11510 8188
rect 11566 8186 11590 8188
rect 11646 8186 11670 8188
rect 11726 8186 11750 8188
rect 11806 8186 11812 8188
rect 11566 8134 11568 8186
rect 11748 8134 11750 8186
rect 11504 8132 11510 8134
rect 11566 8132 11590 8134
rect 11646 8132 11670 8134
rect 11726 8132 11750 8134
rect 11806 8132 11812 8134
rect 11504 8123 11812 8132
rect 11504 7100 11812 7109
rect 11504 7098 11510 7100
rect 11566 7098 11590 7100
rect 11646 7098 11670 7100
rect 11726 7098 11750 7100
rect 11806 7098 11812 7100
rect 11566 7046 11568 7098
rect 11748 7046 11750 7098
rect 11504 7044 11510 7046
rect 11566 7044 11590 7046
rect 11646 7044 11670 7046
rect 11726 7044 11750 7046
rect 11806 7044 11812 7046
rect 11504 7035 11812 7044
rect 11244 6792 11296 6798
rect 11244 6734 11296 6740
rect 10600 6248 10652 6254
rect 10600 6190 10652 6196
rect 9588 6180 9640 6186
rect 9588 6122 9640 6128
rect 9600 5778 9628 6122
rect 9588 5772 9640 5778
rect 9588 5714 9640 5720
rect 10048 5568 10100 5574
rect 10048 5510 10100 5516
rect 10232 5568 10284 5574
rect 10232 5510 10284 5516
rect 9653 5468 9961 5477
rect 9653 5466 9659 5468
rect 9715 5466 9739 5468
rect 9795 5466 9819 5468
rect 9875 5466 9899 5468
rect 9955 5466 9961 5468
rect 9715 5414 9717 5466
rect 9897 5414 9899 5466
rect 9653 5412 9659 5414
rect 9715 5412 9739 5414
rect 9795 5412 9819 5414
rect 9875 5412 9899 5414
rect 9955 5412 9961 5414
rect 9653 5403 9961 5412
rect 10060 5166 10088 5510
rect 9496 5160 9548 5166
rect 9496 5102 9548 5108
rect 10048 5160 10100 5166
rect 10048 5102 10100 5108
rect 10060 4690 10088 5102
rect 10244 4690 10272 5510
rect 11256 5370 11284 6734
rect 11504 6012 11812 6021
rect 11504 6010 11510 6012
rect 11566 6010 11590 6012
rect 11646 6010 11670 6012
rect 11726 6010 11750 6012
rect 11806 6010 11812 6012
rect 11566 5958 11568 6010
rect 11748 5958 11750 6010
rect 11504 5956 11510 5958
rect 11566 5956 11590 5958
rect 11646 5956 11670 5958
rect 11726 5956 11750 5958
rect 11806 5956 11812 5958
rect 11504 5947 11812 5956
rect 11900 5817 11928 13398
rect 12808 13184 12860 13190
rect 12808 13126 12860 13132
rect 11980 12844 12032 12850
rect 11980 12786 12032 12792
rect 11992 11898 12020 12786
rect 12820 12782 12848 13126
rect 12808 12776 12860 12782
rect 12808 12718 12860 12724
rect 12256 12640 12308 12646
rect 12256 12582 12308 12588
rect 12268 12374 12296 12582
rect 12256 12368 12308 12374
rect 12256 12310 12308 12316
rect 12992 12096 13044 12102
rect 12992 12038 13044 12044
rect 11980 11892 12032 11898
rect 11980 11834 12032 11840
rect 12808 11688 12860 11694
rect 12808 11630 12860 11636
rect 12624 11552 12676 11558
rect 12624 11494 12676 11500
rect 12072 11212 12124 11218
rect 12072 11154 12124 11160
rect 11980 10600 12032 10606
rect 11980 10542 12032 10548
rect 11992 10130 12020 10542
rect 12084 10266 12112 11154
rect 12636 11150 12664 11494
rect 12820 11218 12848 11630
rect 12808 11212 12860 11218
rect 12808 11154 12860 11160
rect 13004 11150 13032 12038
rect 12624 11144 12676 11150
rect 12624 11086 12676 11092
rect 12992 11144 13044 11150
rect 12992 11086 13044 11092
rect 12440 10600 12492 10606
rect 12440 10542 12492 10548
rect 12348 10464 12400 10470
rect 12348 10406 12400 10412
rect 12072 10260 12124 10266
rect 12072 10202 12124 10208
rect 12256 10260 12308 10266
rect 12256 10202 12308 10208
rect 11980 10124 12032 10130
rect 11980 10066 12032 10072
rect 12268 9722 12296 10202
rect 12360 10130 12388 10406
rect 12348 10124 12400 10130
rect 12348 10066 12400 10072
rect 12452 9994 12480 10542
rect 12900 10056 12952 10062
rect 12900 9998 12952 10004
rect 12440 9988 12492 9994
rect 12440 9930 12492 9936
rect 12256 9716 12308 9722
rect 12256 9658 12308 9664
rect 12452 9518 12480 9930
rect 12808 9920 12860 9926
rect 12808 9862 12860 9868
rect 12820 9518 12848 9862
rect 12912 9722 12940 9998
rect 12900 9716 12952 9722
rect 12900 9658 12952 9664
rect 12440 9512 12492 9518
rect 12440 9454 12492 9460
rect 12532 9512 12584 9518
rect 12532 9454 12584 9460
rect 12808 9512 12860 9518
rect 12808 9454 12860 9460
rect 12544 9178 12572 9454
rect 12532 9172 12584 9178
rect 12532 9114 12584 9120
rect 12164 9036 12216 9042
rect 12164 8978 12216 8984
rect 12348 9036 12400 9042
rect 12348 8978 12400 8984
rect 12176 8498 12204 8978
rect 12164 8492 12216 8498
rect 12164 8434 12216 8440
rect 12360 8430 12388 8978
rect 12348 8424 12400 8430
rect 12348 8366 12400 8372
rect 12360 7818 12388 8366
rect 12624 8288 12676 8294
rect 12624 8230 12676 8236
rect 12636 7886 12664 8230
rect 12624 7880 12676 7886
rect 12624 7822 12676 7828
rect 12348 7812 12400 7818
rect 12348 7754 12400 7760
rect 12636 7410 12664 7822
rect 12820 7546 12848 9454
rect 13004 9382 13032 11086
rect 13176 9920 13228 9926
rect 13176 9862 13228 9868
rect 12992 9376 13044 9382
rect 12992 9318 13044 9324
rect 13004 9042 13032 9318
rect 13188 9110 13216 9862
rect 13176 9104 13228 9110
rect 13176 9046 13228 9052
rect 12992 9036 13044 9042
rect 12992 8978 13044 8984
rect 13004 7954 13032 8978
rect 13176 8016 13228 8022
rect 13176 7958 13228 7964
rect 12992 7948 13044 7954
rect 12992 7890 13044 7896
rect 13188 7546 13216 7958
rect 12808 7540 12860 7546
rect 12808 7482 12860 7488
rect 13176 7540 13228 7546
rect 13176 7482 13228 7488
rect 13280 7478 13308 15600
rect 13355 15260 13663 15269
rect 13355 15258 13361 15260
rect 13417 15258 13441 15260
rect 13497 15258 13521 15260
rect 13577 15258 13601 15260
rect 13657 15258 13663 15260
rect 13417 15206 13419 15258
rect 13599 15206 13601 15258
rect 13355 15204 13361 15206
rect 13417 15204 13441 15206
rect 13497 15204 13521 15206
rect 13577 15204 13601 15206
rect 13657 15204 13663 15206
rect 13355 15195 13663 15204
rect 15206 14716 15514 14725
rect 15206 14714 15212 14716
rect 15268 14714 15292 14716
rect 15348 14714 15372 14716
rect 15428 14714 15452 14716
rect 15508 14714 15514 14716
rect 15268 14662 15270 14714
rect 15450 14662 15452 14714
rect 15206 14660 15212 14662
rect 15268 14660 15292 14662
rect 15348 14660 15372 14662
rect 15428 14660 15452 14662
rect 15508 14660 15514 14662
rect 15206 14651 15514 14660
rect 15016 14272 15068 14278
rect 15016 14214 15068 14220
rect 13355 14172 13663 14181
rect 13355 14170 13361 14172
rect 13417 14170 13441 14172
rect 13497 14170 13521 14172
rect 13577 14170 13601 14172
rect 13657 14170 13663 14172
rect 13417 14118 13419 14170
rect 13599 14118 13601 14170
rect 13355 14116 13361 14118
rect 13417 14116 13441 14118
rect 13497 14116 13521 14118
rect 13577 14116 13601 14118
rect 13657 14116 13663 14118
rect 13355 14107 13663 14116
rect 15028 13977 15056 14214
rect 15014 13968 15070 13977
rect 15014 13903 15070 13912
rect 15206 13628 15514 13637
rect 15206 13626 15212 13628
rect 15268 13626 15292 13628
rect 15348 13626 15372 13628
rect 15428 13626 15452 13628
rect 15508 13626 15514 13628
rect 15268 13574 15270 13626
rect 15450 13574 15452 13626
rect 15206 13572 15212 13574
rect 15268 13572 15292 13574
rect 15348 13572 15372 13574
rect 15428 13572 15452 13574
rect 15508 13572 15514 13574
rect 15206 13563 15514 13572
rect 15016 13184 15068 13190
rect 15014 13152 15016 13161
rect 15068 13152 15070 13161
rect 13355 13084 13663 13093
rect 15014 13087 15070 13096
rect 13355 13082 13361 13084
rect 13417 13082 13441 13084
rect 13497 13082 13521 13084
rect 13577 13082 13601 13084
rect 13657 13082 13663 13084
rect 13417 13030 13419 13082
rect 13599 13030 13601 13082
rect 13355 13028 13361 13030
rect 13417 13028 13441 13030
rect 13497 13028 13521 13030
rect 13577 13028 13601 13030
rect 13657 13028 13663 13030
rect 13355 13019 13663 13028
rect 15016 12776 15068 12782
rect 15016 12718 15068 12724
rect 14740 12708 14792 12714
rect 14740 12650 14792 12656
rect 14752 12238 14780 12650
rect 15028 12345 15056 12718
rect 15206 12540 15514 12549
rect 15206 12538 15212 12540
rect 15268 12538 15292 12540
rect 15348 12538 15372 12540
rect 15428 12538 15452 12540
rect 15508 12538 15514 12540
rect 15268 12486 15270 12538
rect 15450 12486 15452 12538
rect 15206 12484 15212 12486
rect 15268 12484 15292 12486
rect 15348 12484 15372 12486
rect 15428 12484 15452 12486
rect 15508 12484 15514 12486
rect 15206 12475 15514 12484
rect 15014 12336 15070 12345
rect 15014 12271 15070 12280
rect 13728 12232 13780 12238
rect 13728 12174 13780 12180
rect 14740 12232 14792 12238
rect 14740 12174 14792 12180
rect 13355 11996 13663 12005
rect 13355 11994 13361 11996
rect 13417 11994 13441 11996
rect 13497 11994 13521 11996
rect 13577 11994 13601 11996
rect 13657 11994 13663 11996
rect 13417 11942 13419 11994
rect 13599 11942 13601 11994
rect 13355 11940 13361 11942
rect 13417 11940 13441 11942
rect 13497 11940 13521 11942
rect 13577 11940 13601 11942
rect 13657 11940 13663 11942
rect 13355 11931 13663 11940
rect 13740 11286 13768 12174
rect 13728 11280 13780 11286
rect 13728 11222 13780 11228
rect 13355 10908 13663 10917
rect 13355 10906 13361 10908
rect 13417 10906 13441 10908
rect 13497 10906 13521 10908
rect 13577 10906 13601 10908
rect 13657 10906 13663 10908
rect 13417 10854 13419 10906
rect 13599 10854 13601 10906
rect 13355 10852 13361 10854
rect 13417 10852 13441 10854
rect 13497 10852 13521 10854
rect 13577 10852 13601 10854
rect 13657 10852 13663 10854
rect 13355 10843 13663 10852
rect 13355 9820 13663 9829
rect 13355 9818 13361 9820
rect 13417 9818 13441 9820
rect 13497 9818 13521 9820
rect 13577 9818 13601 9820
rect 13657 9818 13663 9820
rect 13417 9766 13419 9818
rect 13599 9766 13601 9818
rect 13355 9764 13361 9766
rect 13417 9764 13441 9766
rect 13497 9764 13521 9766
rect 13577 9764 13601 9766
rect 13657 9764 13663 9766
rect 13355 9755 13663 9764
rect 13740 9110 13768 11222
rect 13728 9104 13780 9110
rect 13728 9046 13780 9052
rect 13355 8732 13663 8741
rect 13355 8730 13361 8732
rect 13417 8730 13441 8732
rect 13497 8730 13521 8732
rect 13577 8730 13601 8732
rect 13657 8730 13663 8732
rect 13417 8678 13419 8730
rect 13599 8678 13601 8730
rect 13355 8676 13361 8678
rect 13417 8676 13441 8678
rect 13497 8676 13521 8678
rect 13577 8676 13601 8678
rect 13657 8676 13663 8678
rect 13355 8667 13663 8676
rect 13740 8022 13768 9046
rect 13728 8016 13780 8022
rect 13726 7984 13728 7993
rect 13780 7984 13782 7993
rect 13726 7919 13782 7928
rect 13355 7644 13663 7653
rect 13355 7642 13361 7644
rect 13417 7642 13441 7644
rect 13497 7642 13521 7644
rect 13577 7642 13601 7644
rect 13657 7642 13663 7644
rect 13417 7590 13419 7642
rect 13599 7590 13601 7642
rect 13355 7588 13361 7590
rect 13417 7588 13441 7590
rect 13497 7588 13521 7590
rect 13577 7588 13601 7590
rect 13657 7588 13663 7590
rect 13355 7579 13663 7588
rect 13268 7472 13320 7478
rect 14752 7449 14780 12174
rect 15660 11824 15712 11830
rect 15660 11766 15712 11772
rect 15672 11529 15700 11766
rect 15658 11520 15714 11529
rect 15206 11452 15514 11461
rect 15658 11455 15714 11464
rect 15206 11450 15212 11452
rect 15268 11450 15292 11452
rect 15348 11450 15372 11452
rect 15428 11450 15452 11452
rect 15508 11450 15514 11452
rect 15268 11398 15270 11450
rect 15450 11398 15452 11450
rect 15206 11396 15212 11398
rect 15268 11396 15292 11398
rect 15348 11396 15372 11398
rect 15428 11396 15452 11398
rect 15508 11396 15514 11398
rect 15206 11387 15514 11396
rect 14924 11144 14976 11150
rect 14924 11086 14976 11092
rect 13268 7414 13320 7420
rect 14738 7440 14794 7449
rect 12624 7404 12676 7410
rect 14738 7375 14794 7384
rect 12624 7346 12676 7352
rect 12808 7336 12860 7342
rect 12808 7278 12860 7284
rect 13268 7336 13320 7342
rect 13268 7278 13320 7284
rect 13820 7336 13872 7342
rect 13820 7278 13872 7284
rect 12820 6866 12848 7278
rect 12900 7268 12952 7274
rect 12900 7210 12952 7216
rect 11980 6860 12032 6866
rect 11980 6802 12032 6808
rect 12808 6860 12860 6866
rect 12808 6802 12860 6808
rect 11992 6730 12020 6802
rect 11980 6724 12032 6730
rect 11980 6666 12032 6672
rect 11886 5808 11942 5817
rect 11886 5743 11942 5752
rect 11992 5642 12020 6666
rect 12912 6254 12940 7210
rect 13280 6662 13308 7278
rect 13728 7200 13780 7206
rect 13728 7142 13780 7148
rect 13268 6656 13320 6662
rect 13268 6598 13320 6604
rect 13355 6556 13663 6565
rect 13355 6554 13361 6556
rect 13417 6554 13441 6556
rect 13497 6554 13521 6556
rect 13577 6554 13601 6556
rect 13657 6554 13663 6556
rect 13417 6502 13419 6554
rect 13599 6502 13601 6554
rect 13355 6500 13361 6502
rect 13417 6500 13441 6502
rect 13497 6500 13521 6502
rect 13577 6500 13601 6502
rect 13657 6500 13663 6502
rect 13355 6491 13663 6500
rect 13740 6254 13768 7142
rect 12900 6248 12952 6254
rect 12900 6190 12952 6196
rect 13728 6248 13780 6254
rect 13728 6190 13780 6196
rect 13544 6112 13596 6118
rect 13544 6054 13596 6060
rect 13556 5846 13584 6054
rect 13544 5840 13596 5846
rect 13544 5782 13596 5788
rect 12992 5704 13044 5710
rect 12992 5646 13044 5652
rect 11980 5636 12032 5642
rect 11980 5578 12032 5584
rect 11244 5364 11296 5370
rect 11244 5306 11296 5312
rect 13004 5302 13032 5646
rect 13355 5468 13663 5477
rect 13355 5466 13361 5468
rect 13417 5466 13441 5468
rect 13497 5466 13521 5468
rect 13577 5466 13601 5468
rect 13657 5466 13663 5468
rect 13417 5414 13419 5466
rect 13599 5414 13601 5466
rect 13355 5412 13361 5414
rect 13417 5412 13441 5414
rect 13497 5412 13521 5414
rect 13577 5412 13601 5414
rect 13657 5412 13663 5414
rect 13355 5403 13663 5412
rect 13740 5370 13768 6190
rect 13832 6186 13860 7278
rect 13912 6656 13964 6662
rect 14936 6633 14964 11086
rect 15014 10704 15070 10713
rect 15014 10639 15016 10648
rect 15068 10639 15070 10648
rect 15016 10610 15068 10616
rect 15206 10364 15514 10373
rect 15206 10362 15212 10364
rect 15268 10362 15292 10364
rect 15348 10362 15372 10364
rect 15428 10362 15452 10364
rect 15508 10362 15514 10364
rect 15268 10310 15270 10362
rect 15450 10310 15452 10362
rect 15206 10308 15212 10310
rect 15268 10308 15292 10310
rect 15348 10308 15372 10310
rect 15428 10308 15452 10310
rect 15508 10308 15514 10310
rect 15206 10299 15514 10308
rect 15016 9920 15068 9926
rect 15014 9888 15016 9897
rect 15068 9888 15070 9897
rect 15014 9823 15070 9832
rect 15016 9512 15068 9518
rect 15016 9454 15068 9460
rect 15028 9081 15056 9454
rect 15206 9276 15514 9285
rect 15206 9274 15212 9276
rect 15268 9274 15292 9276
rect 15348 9274 15372 9276
rect 15428 9274 15452 9276
rect 15508 9274 15514 9276
rect 15268 9222 15270 9274
rect 15450 9222 15452 9274
rect 15206 9220 15212 9222
rect 15268 9220 15292 9222
rect 15348 9220 15372 9222
rect 15428 9220 15452 9222
rect 15508 9220 15514 9222
rect 15206 9211 15514 9220
rect 15014 9072 15070 9081
rect 15014 9007 15070 9016
rect 15568 8968 15620 8974
rect 15568 8910 15620 8916
rect 15206 8188 15514 8197
rect 15206 8186 15212 8188
rect 15268 8186 15292 8188
rect 15348 8186 15372 8188
rect 15428 8186 15452 8188
rect 15508 8186 15514 8188
rect 15268 8134 15270 8186
rect 15450 8134 15452 8186
rect 15206 8132 15212 8134
rect 15268 8132 15292 8134
rect 15348 8132 15372 8134
rect 15428 8132 15452 8134
rect 15508 8132 15514 8134
rect 15206 8123 15514 8132
rect 15016 8016 15068 8022
rect 15016 7958 15068 7964
rect 15028 6905 15056 7958
rect 15206 7100 15514 7109
rect 15206 7098 15212 7100
rect 15268 7098 15292 7100
rect 15348 7098 15372 7100
rect 15428 7098 15452 7100
rect 15508 7098 15514 7100
rect 15268 7046 15270 7098
rect 15450 7046 15452 7098
rect 15206 7044 15212 7046
rect 15268 7044 15292 7046
rect 15348 7044 15372 7046
rect 15428 7044 15452 7046
rect 15508 7044 15514 7046
rect 15206 7035 15514 7044
rect 15014 6896 15070 6905
rect 15014 6831 15070 6840
rect 13912 6598 13964 6604
rect 14922 6624 14978 6633
rect 13924 6254 13952 6598
rect 14922 6559 14978 6568
rect 13912 6248 13964 6254
rect 13912 6190 13964 6196
rect 13820 6180 13872 6186
rect 13820 6122 13872 6128
rect 13728 5364 13780 5370
rect 13728 5306 13780 5312
rect 12992 5296 13044 5302
rect 12992 5238 13044 5244
rect 11336 5160 11388 5166
rect 11336 5102 11388 5108
rect 11428 5160 11480 5166
rect 11428 5102 11480 5108
rect 12164 5160 12216 5166
rect 12164 5102 12216 5108
rect 12808 5160 12860 5166
rect 12808 5102 12860 5108
rect 11060 5092 11112 5098
rect 11060 5034 11112 5040
rect 10692 5024 10744 5030
rect 10692 4966 10744 4972
rect 10704 4826 10732 4966
rect 10692 4820 10744 4826
rect 10692 4762 10744 4768
rect 10048 4684 10100 4690
rect 10048 4626 10100 4632
rect 10232 4684 10284 4690
rect 10232 4626 10284 4632
rect 11072 4622 11100 5034
rect 11348 4826 11376 5102
rect 11336 4820 11388 4826
rect 11336 4762 11388 4768
rect 11440 4690 11468 5102
rect 11504 4924 11812 4933
rect 11504 4922 11510 4924
rect 11566 4922 11590 4924
rect 11646 4922 11670 4924
rect 11726 4922 11750 4924
rect 11806 4922 11812 4924
rect 11566 4870 11568 4922
rect 11748 4870 11750 4922
rect 11504 4868 11510 4870
rect 11566 4868 11590 4870
rect 11646 4868 11670 4870
rect 11726 4868 11750 4870
rect 11806 4868 11812 4870
rect 11504 4859 11812 4868
rect 11244 4684 11296 4690
rect 11244 4626 11296 4632
rect 11336 4684 11388 4690
rect 11336 4626 11388 4632
rect 11428 4684 11480 4690
rect 11428 4626 11480 4632
rect 11520 4684 11572 4690
rect 11520 4626 11572 4632
rect 11060 4616 11112 4622
rect 11060 4558 11112 4564
rect 10508 4480 10560 4486
rect 10508 4422 10560 4428
rect 9653 4380 9961 4389
rect 9653 4378 9659 4380
rect 9715 4378 9739 4380
rect 9795 4378 9819 4380
rect 9875 4378 9899 4380
rect 9955 4378 9961 4380
rect 9715 4326 9717 4378
rect 9897 4326 9899 4378
rect 9653 4324 9659 4326
rect 9715 4324 9739 4326
rect 9795 4324 9819 4326
rect 9875 4324 9899 4326
rect 9955 4324 9961 4326
rect 9653 4315 9961 4324
rect 10520 4214 10548 4422
rect 11256 4214 11284 4626
rect 10508 4208 10560 4214
rect 10508 4150 10560 4156
rect 11244 4208 11296 4214
rect 11244 4150 11296 4156
rect 10232 4004 10284 4010
rect 10232 3946 10284 3952
rect 9680 3936 9732 3942
rect 9680 3878 9732 3884
rect 10244 3890 10272 3946
rect 10520 3942 10548 4150
rect 11256 4078 11284 4150
rect 11244 4072 11296 4078
rect 11244 4014 11296 4020
rect 10508 3936 10560 3942
rect 9692 3738 9720 3878
rect 10244 3862 10364 3890
rect 10508 3878 10560 3884
rect 9680 3732 9732 3738
rect 9680 3674 9732 3680
rect 8576 3596 8628 3602
rect 8576 3538 8628 3544
rect 9036 3596 9088 3602
rect 9036 3538 9088 3544
rect 9128 3596 9180 3602
rect 9128 3538 9180 3544
rect 9312 3596 9364 3602
rect 9312 3538 9364 3544
rect 6644 2916 6696 2922
rect 6644 2858 6696 2864
rect 7656 2916 7708 2922
rect 7656 2858 7708 2864
rect 4100 2748 4408 2757
rect 4100 2746 4106 2748
rect 4162 2746 4186 2748
rect 4242 2746 4266 2748
rect 4322 2746 4346 2748
rect 4402 2746 4408 2748
rect 4162 2694 4164 2746
rect 4344 2694 4346 2746
rect 4100 2692 4106 2694
rect 4162 2692 4186 2694
rect 4242 2692 4266 2694
rect 4322 2692 4346 2694
rect 4402 2692 4408 2694
rect 4100 2683 4408 2692
rect 6656 2650 6684 2858
rect 8208 2848 8260 2854
rect 8208 2790 8260 2796
rect 7802 2748 8110 2757
rect 7802 2746 7808 2748
rect 7864 2746 7888 2748
rect 7944 2746 7968 2748
rect 8024 2746 8048 2748
rect 8104 2746 8110 2748
rect 7864 2694 7866 2746
rect 8046 2694 8048 2746
rect 7802 2692 7808 2694
rect 7864 2692 7888 2694
rect 7944 2692 7968 2694
rect 8024 2692 8048 2694
rect 8104 2692 8110 2694
rect 7802 2683 8110 2692
rect 6644 2644 6696 2650
rect 6644 2586 6696 2592
rect 8220 2582 8248 2790
rect 8208 2576 8260 2582
rect 8208 2518 8260 2524
rect 8298 2544 8354 2553
rect 8298 2479 8300 2488
rect 8352 2479 8354 2488
rect 8300 2450 8352 2456
rect 2249 2204 2557 2213
rect 2249 2202 2255 2204
rect 2311 2202 2335 2204
rect 2391 2202 2415 2204
rect 2471 2202 2495 2204
rect 2551 2202 2557 2204
rect 2311 2150 2313 2202
rect 2493 2150 2495 2202
rect 2249 2148 2255 2150
rect 2311 2148 2335 2150
rect 2391 2148 2415 2150
rect 2471 2148 2495 2150
rect 2551 2148 2557 2150
rect 2249 2139 2557 2148
rect 5951 2204 6259 2213
rect 5951 2202 5957 2204
rect 6013 2202 6037 2204
rect 6093 2202 6117 2204
rect 6173 2202 6197 2204
rect 6253 2202 6259 2204
rect 6013 2150 6015 2202
rect 6195 2150 6197 2202
rect 5951 2148 5957 2150
rect 6013 2148 6037 2150
rect 6093 2148 6117 2150
rect 6173 2148 6197 2150
rect 6253 2148 6259 2150
rect 5951 2139 6259 2148
rect 8312 1902 8340 2450
rect 8300 1896 8352 1902
rect 8300 1838 8352 1844
rect 7656 1760 7708 1766
rect 7656 1702 7708 1708
rect 4100 1660 4408 1669
rect 4100 1658 4106 1660
rect 4162 1658 4186 1660
rect 4242 1658 4266 1660
rect 4322 1658 4346 1660
rect 4402 1658 4408 1660
rect 4162 1606 4164 1658
rect 4344 1606 4346 1658
rect 4100 1604 4106 1606
rect 4162 1604 4186 1606
rect 4242 1604 4266 1606
rect 4322 1604 4346 1606
rect 4402 1604 4408 1606
rect 4100 1595 4408 1604
rect 7196 1352 7248 1358
rect 7196 1294 7248 1300
rect 2249 1116 2557 1125
rect 2249 1114 2255 1116
rect 2311 1114 2335 1116
rect 2391 1114 2415 1116
rect 2471 1114 2495 1116
rect 2551 1114 2557 1116
rect 2311 1062 2313 1114
rect 2493 1062 2495 1114
rect 2249 1060 2255 1062
rect 2311 1060 2335 1062
rect 2391 1060 2415 1062
rect 2471 1060 2495 1062
rect 2551 1060 2557 1062
rect 2249 1051 2557 1060
rect 5951 1116 6259 1125
rect 5951 1114 5957 1116
rect 6013 1114 6037 1116
rect 6093 1114 6117 1116
rect 6173 1114 6197 1116
rect 6253 1114 6259 1116
rect 6013 1062 6015 1114
rect 6195 1062 6197 1114
rect 5951 1060 5957 1062
rect 6013 1060 6037 1062
rect 6093 1060 6117 1062
rect 6173 1060 6197 1062
rect 6253 1060 6259 1062
rect 5951 1051 6259 1060
rect 7208 1018 7236 1294
rect 7196 1012 7248 1018
rect 7196 954 7248 960
rect 7668 814 7696 1702
rect 7802 1660 8110 1669
rect 7802 1658 7808 1660
rect 7864 1658 7888 1660
rect 7944 1658 7968 1660
rect 8024 1658 8048 1660
rect 8104 1658 8110 1660
rect 7864 1606 7866 1658
rect 8046 1606 8048 1658
rect 7802 1604 7808 1606
rect 7864 1604 7888 1606
rect 7944 1604 7968 1606
rect 8024 1604 8048 1606
rect 8104 1604 8110 1606
rect 7802 1595 8110 1604
rect 8588 1018 8616 3538
rect 8760 2508 8812 2514
rect 8760 2450 8812 2456
rect 8772 1426 8800 2450
rect 9140 2310 9168 3538
rect 9653 3292 9961 3301
rect 9653 3290 9659 3292
rect 9715 3290 9739 3292
rect 9795 3290 9819 3292
rect 9875 3290 9899 3292
rect 9955 3290 9961 3292
rect 9715 3238 9717 3290
rect 9897 3238 9899 3290
rect 9653 3236 9659 3238
rect 9715 3236 9739 3238
rect 9795 3236 9819 3238
rect 9875 3236 9899 3238
rect 9955 3236 9961 3238
rect 9653 3227 9961 3236
rect 9496 2984 9548 2990
rect 9496 2926 9548 2932
rect 9312 2848 9364 2854
rect 9312 2790 9364 2796
rect 9324 2514 9352 2790
rect 9312 2508 9364 2514
rect 9312 2450 9364 2456
rect 9128 2304 9180 2310
rect 9128 2246 9180 2252
rect 9140 1970 9168 2246
rect 9508 2106 9536 2926
rect 10336 2582 10364 3862
rect 11348 3602 11376 4626
rect 11440 3942 11468 4626
rect 11532 4214 11560 4626
rect 12176 4554 12204 5102
rect 12820 4758 12848 5102
rect 12808 4752 12860 4758
rect 12808 4694 12860 4700
rect 12164 4548 12216 4554
rect 12164 4490 12216 4496
rect 11520 4208 11572 4214
rect 11520 4150 11572 4156
rect 12808 4004 12860 4010
rect 12808 3946 12860 3952
rect 11428 3936 11480 3942
rect 11428 3878 11480 3884
rect 11336 3596 11388 3602
rect 11336 3538 11388 3544
rect 10324 2576 10376 2582
rect 10324 2518 10376 2524
rect 10140 2304 10192 2310
rect 10140 2246 10192 2252
rect 9653 2204 9961 2213
rect 9653 2202 9659 2204
rect 9715 2202 9739 2204
rect 9795 2202 9819 2204
rect 9875 2202 9899 2204
rect 9955 2202 9961 2204
rect 9715 2150 9717 2202
rect 9897 2150 9899 2202
rect 9653 2148 9659 2150
rect 9715 2148 9739 2150
rect 9795 2148 9819 2150
rect 9875 2148 9899 2150
rect 9955 2148 9961 2150
rect 9653 2139 9961 2148
rect 9496 2100 9548 2106
rect 9496 2042 9548 2048
rect 10152 1970 10180 2246
rect 8852 1964 8904 1970
rect 8852 1906 8904 1912
rect 9128 1964 9180 1970
rect 9128 1906 9180 1912
rect 10140 1964 10192 1970
rect 10140 1906 10192 1912
rect 8864 1562 8892 1906
rect 9140 1766 9168 1906
rect 10046 1864 10102 1873
rect 10046 1799 10048 1808
rect 10100 1799 10102 1808
rect 10048 1770 10100 1776
rect 9128 1760 9180 1766
rect 9128 1702 9180 1708
rect 8852 1556 8904 1562
rect 8852 1498 8904 1504
rect 8760 1420 8812 1426
rect 8760 1362 8812 1368
rect 9036 1352 9088 1358
rect 9036 1294 9088 1300
rect 9048 1018 9076 1294
rect 9653 1116 9961 1125
rect 9653 1114 9659 1116
rect 9715 1114 9739 1116
rect 9795 1114 9819 1116
rect 9875 1114 9899 1116
rect 9955 1114 9961 1116
rect 9715 1062 9717 1114
rect 9897 1062 9899 1114
rect 9653 1060 9659 1062
rect 9715 1060 9739 1062
rect 9795 1060 9819 1062
rect 9875 1060 9899 1062
rect 9955 1060 9961 1062
rect 9653 1051 9961 1060
rect 8576 1012 8628 1018
rect 8576 954 8628 960
rect 9036 1012 9088 1018
rect 9036 954 9088 960
rect 10060 882 10088 1770
rect 10140 1760 10192 1766
rect 10140 1702 10192 1708
rect 10152 882 10180 1702
rect 10336 1494 10364 2518
rect 10876 2440 10928 2446
rect 10876 2382 10928 2388
rect 10888 1834 10916 2382
rect 11348 2106 11376 3538
rect 11440 3534 11468 3878
rect 11504 3836 11812 3845
rect 11504 3834 11510 3836
rect 11566 3834 11590 3836
rect 11646 3834 11670 3836
rect 11726 3834 11750 3836
rect 11806 3834 11812 3836
rect 11566 3782 11568 3834
rect 11748 3782 11750 3834
rect 11504 3780 11510 3782
rect 11566 3780 11590 3782
rect 11646 3780 11670 3782
rect 11726 3780 11750 3782
rect 11806 3780 11812 3782
rect 11504 3771 11812 3780
rect 12820 3738 12848 3946
rect 12808 3732 12860 3738
rect 12808 3674 12860 3680
rect 13004 3602 13032 5238
rect 13728 5160 13780 5166
rect 13728 5102 13780 5108
rect 13176 5024 13228 5030
rect 13176 4966 13228 4972
rect 13084 4276 13136 4282
rect 13084 4218 13136 4224
rect 13096 4185 13124 4218
rect 13082 4176 13138 4185
rect 13188 4146 13216 4966
rect 13740 4690 13768 5102
rect 13728 4684 13780 4690
rect 13728 4626 13780 4632
rect 13268 4480 13320 4486
rect 13268 4422 13320 4428
rect 13082 4111 13138 4120
rect 13176 4140 13228 4146
rect 13176 4082 13228 4088
rect 13280 3670 13308 4422
rect 13355 4380 13663 4389
rect 13355 4378 13361 4380
rect 13417 4378 13441 4380
rect 13497 4378 13521 4380
rect 13577 4378 13601 4380
rect 13657 4378 13663 4380
rect 13417 4326 13419 4378
rect 13599 4326 13601 4378
rect 13355 4324 13361 4326
rect 13417 4324 13441 4326
rect 13497 4324 13521 4326
rect 13577 4324 13601 4326
rect 13657 4324 13663 4326
rect 13355 4315 13663 4324
rect 13728 4208 13780 4214
rect 13728 4154 13780 4156
rect 13832 4154 13860 6122
rect 15206 6012 15514 6021
rect 15206 6010 15212 6012
rect 15268 6010 15292 6012
rect 15348 6010 15372 6012
rect 15428 6010 15452 6012
rect 15508 6010 15514 6012
rect 15268 5958 15270 6010
rect 15450 5958 15452 6010
rect 15206 5956 15212 5958
rect 15268 5956 15292 5958
rect 15348 5956 15372 5958
rect 15428 5956 15452 5958
rect 15508 5956 15514 5958
rect 15206 5947 15514 5956
rect 15016 5908 15068 5914
rect 15016 5850 15068 5856
rect 13912 5840 13964 5846
rect 13910 5808 13912 5817
rect 13964 5808 13966 5817
rect 13966 5766 14044 5794
rect 13910 5743 13966 5752
rect 13912 4684 13964 4690
rect 13912 4626 13964 4632
rect 13924 4282 13952 4626
rect 13912 4276 13964 4282
rect 13912 4218 13964 4224
rect 13728 4150 13860 4154
rect 13740 4126 13860 4150
rect 13832 4010 13860 4126
rect 13910 4176 13966 4185
rect 13910 4111 13966 4120
rect 13924 4078 13952 4111
rect 13912 4072 13964 4078
rect 13912 4014 13964 4020
rect 13820 4004 13872 4010
rect 13820 3946 13872 3952
rect 13268 3664 13320 3670
rect 13268 3606 13320 3612
rect 12348 3596 12400 3602
rect 12348 3538 12400 3544
rect 12992 3596 13044 3602
rect 12992 3538 13044 3544
rect 11428 3528 11480 3534
rect 11428 3470 11480 3476
rect 12360 3058 12388 3538
rect 12440 3528 12492 3534
rect 12440 3470 12492 3476
rect 12348 3052 12400 3058
rect 12348 2994 12400 3000
rect 12452 2990 12480 3470
rect 12440 2984 12492 2990
rect 12440 2926 12492 2932
rect 11504 2748 11812 2757
rect 11504 2746 11510 2748
rect 11566 2746 11590 2748
rect 11646 2746 11670 2748
rect 11726 2746 11750 2748
rect 11806 2746 11812 2748
rect 11566 2694 11568 2746
rect 11748 2694 11750 2746
rect 11504 2692 11510 2694
rect 11566 2692 11590 2694
rect 11646 2692 11670 2694
rect 11726 2692 11750 2694
rect 11806 2692 11812 2694
rect 11504 2683 11812 2692
rect 11428 2304 11480 2310
rect 11428 2246 11480 2252
rect 11336 2100 11388 2106
rect 11336 2042 11388 2048
rect 11152 2032 11204 2038
rect 11152 1974 11204 1980
rect 10876 1828 10928 1834
rect 10876 1770 10928 1776
rect 10324 1488 10376 1494
rect 10324 1430 10376 1436
rect 10888 1426 10916 1770
rect 10876 1420 10928 1426
rect 10876 1362 10928 1368
rect 11164 1358 11192 1974
rect 11152 1352 11204 1358
rect 11152 1294 11204 1300
rect 10508 1216 10560 1222
rect 10508 1158 10560 1164
rect 10048 876 10100 882
rect 10048 818 10100 824
rect 10140 876 10192 882
rect 10140 818 10192 824
rect 10520 814 10548 1158
rect 11440 814 11468 2246
rect 12072 1896 12124 1902
rect 12072 1838 12124 1844
rect 12348 1896 12400 1902
rect 12348 1838 12400 1844
rect 11504 1660 11812 1669
rect 11504 1658 11510 1660
rect 11566 1658 11590 1660
rect 11646 1658 11670 1660
rect 11726 1658 11750 1660
rect 11806 1658 11812 1660
rect 11566 1606 11568 1658
rect 11748 1606 11750 1658
rect 11504 1604 11510 1606
rect 11566 1604 11590 1606
rect 11646 1604 11670 1606
rect 11726 1604 11750 1606
rect 11806 1604 11812 1606
rect 11504 1595 11812 1604
rect 12084 1018 12112 1838
rect 12360 1766 12388 1838
rect 12348 1760 12400 1766
rect 12348 1702 12400 1708
rect 12360 1562 12388 1702
rect 12348 1556 12400 1562
rect 12348 1498 12400 1504
rect 12164 1352 12216 1358
rect 12164 1294 12216 1300
rect 12072 1012 12124 1018
rect 12072 954 12124 960
rect 12176 814 12204 1294
rect 12360 950 12388 1498
rect 12452 1426 12480 2926
rect 12716 2848 12768 2854
rect 12716 2790 12768 2796
rect 12728 2514 12756 2790
rect 13004 2650 13032 3538
rect 13355 3292 13663 3301
rect 13355 3290 13361 3292
rect 13417 3290 13441 3292
rect 13497 3290 13521 3292
rect 13577 3290 13601 3292
rect 13657 3290 13663 3292
rect 13417 3238 13419 3290
rect 13599 3238 13601 3290
rect 13355 3236 13361 3238
rect 13417 3236 13441 3238
rect 13497 3236 13521 3238
rect 13577 3236 13601 3238
rect 13657 3236 13663 3238
rect 13355 3227 13663 3236
rect 12992 2644 13044 2650
rect 12992 2586 13044 2592
rect 13004 2514 13032 2586
rect 12716 2508 12768 2514
rect 12716 2450 12768 2456
rect 12992 2508 13044 2514
rect 12992 2450 13044 2456
rect 12532 2440 12584 2446
rect 12532 2382 12584 2388
rect 12544 1970 12572 2382
rect 12532 1964 12584 1970
rect 12532 1906 12584 1912
rect 12624 1828 12676 1834
rect 12624 1770 12676 1776
rect 12440 1420 12492 1426
rect 12440 1362 12492 1368
rect 12636 1018 12664 1770
rect 12728 1766 12756 2450
rect 12900 2304 12952 2310
rect 12900 2246 12952 2252
rect 12912 1970 12940 2246
rect 12900 1964 12952 1970
rect 12900 1906 12952 1912
rect 12716 1760 12768 1766
rect 12716 1702 12768 1708
rect 12808 1760 12860 1766
rect 12808 1702 12860 1708
rect 12716 1216 12768 1222
rect 12716 1158 12768 1164
rect 12624 1012 12676 1018
rect 12624 954 12676 960
rect 12348 944 12400 950
rect 12348 886 12400 892
rect 12728 882 12756 1158
rect 12820 1018 12848 1702
rect 13004 1426 13032 2450
rect 13268 2440 13320 2446
rect 13268 2382 13320 2388
rect 13280 2106 13308 2382
rect 13355 2204 13663 2213
rect 13355 2202 13361 2204
rect 13417 2202 13441 2204
rect 13497 2202 13521 2204
rect 13577 2202 13601 2204
rect 13657 2202 13663 2204
rect 13417 2150 13419 2202
rect 13599 2150 13601 2202
rect 13355 2148 13361 2150
rect 13417 2148 13441 2150
rect 13497 2148 13521 2150
rect 13577 2148 13601 2150
rect 13657 2148 13663 2150
rect 13355 2139 13663 2148
rect 13268 2100 13320 2106
rect 13268 2042 13320 2048
rect 13924 1902 13952 4014
rect 14016 3670 14044 5766
rect 15028 5710 15056 5850
rect 15580 5817 15608 8910
rect 15660 8424 15712 8430
rect 15660 8366 15712 8372
rect 15672 8265 15700 8366
rect 15658 8256 15714 8265
rect 15658 8191 15714 8200
rect 15934 6896 15990 6905
rect 15934 6831 15990 6840
rect 15566 5808 15622 5817
rect 15566 5743 15622 5752
rect 15016 5704 15068 5710
rect 15016 5646 15068 5652
rect 15028 4185 15056 5646
rect 15948 5001 15976 6831
rect 15934 4992 15990 5001
rect 15206 4924 15514 4933
rect 15934 4927 15990 4936
rect 15206 4922 15212 4924
rect 15268 4922 15292 4924
rect 15348 4922 15372 4924
rect 15428 4922 15452 4924
rect 15508 4922 15514 4924
rect 15268 4870 15270 4922
rect 15450 4870 15452 4922
rect 15206 4868 15212 4870
rect 15268 4868 15292 4870
rect 15348 4868 15372 4870
rect 15428 4868 15452 4870
rect 15508 4868 15514 4870
rect 15206 4859 15514 4868
rect 15014 4176 15070 4185
rect 15014 4111 15070 4120
rect 15206 3836 15514 3845
rect 15206 3834 15212 3836
rect 15268 3834 15292 3836
rect 15348 3834 15372 3836
rect 15428 3834 15452 3836
rect 15508 3834 15514 3836
rect 15268 3782 15270 3834
rect 15450 3782 15452 3834
rect 15206 3780 15212 3782
rect 15268 3780 15292 3782
rect 15348 3780 15372 3782
rect 15428 3780 15452 3782
rect 15508 3780 15514 3782
rect 15206 3771 15514 3780
rect 14004 3664 14056 3670
rect 14004 3606 14056 3612
rect 14016 2582 14044 3606
rect 15016 3528 15068 3534
rect 15016 3470 15068 3476
rect 15028 3369 15056 3470
rect 15014 3360 15070 3369
rect 15014 3295 15070 3304
rect 15206 2748 15514 2757
rect 15206 2746 15212 2748
rect 15268 2746 15292 2748
rect 15348 2746 15372 2748
rect 15428 2746 15452 2748
rect 15508 2746 15514 2748
rect 15268 2694 15270 2746
rect 15450 2694 15452 2746
rect 15206 2692 15212 2694
rect 15268 2692 15292 2694
rect 15348 2692 15372 2694
rect 15428 2692 15452 2694
rect 15508 2692 15514 2694
rect 15206 2683 15514 2692
rect 14004 2576 14056 2582
rect 14004 2518 14056 2524
rect 15014 2544 15070 2553
rect 15014 2479 15016 2488
rect 15068 2479 15070 2488
rect 15016 2450 15068 2456
rect 13084 1896 13136 1902
rect 13084 1838 13136 1844
rect 13912 1896 13964 1902
rect 13912 1838 13964 1844
rect 15014 1864 15070 1873
rect 12992 1420 13044 1426
rect 12992 1362 13044 1368
rect 12808 1012 12860 1018
rect 12808 954 12860 960
rect 12716 876 12768 882
rect 12716 818 12768 824
rect 13096 814 13124 1838
rect 15014 1799 15070 1808
rect 15028 1494 15056 1799
rect 15658 1728 15714 1737
rect 15206 1660 15514 1669
rect 15658 1663 15714 1672
rect 15206 1658 15212 1660
rect 15268 1658 15292 1660
rect 15348 1658 15372 1660
rect 15428 1658 15452 1660
rect 15508 1658 15514 1660
rect 15268 1606 15270 1658
rect 15450 1606 15452 1658
rect 15206 1604 15212 1606
rect 15268 1604 15292 1606
rect 15348 1604 15372 1606
rect 15428 1604 15452 1606
rect 15508 1604 15514 1606
rect 15206 1595 15514 1604
rect 15672 1494 15700 1663
rect 15016 1488 15068 1494
rect 15016 1430 15068 1436
rect 15660 1488 15712 1494
rect 15660 1430 15712 1436
rect 13268 1352 13320 1358
rect 13268 1294 13320 1300
rect 13280 1018 13308 1294
rect 13355 1116 13663 1125
rect 13355 1114 13361 1116
rect 13417 1114 13441 1116
rect 13497 1114 13521 1116
rect 13577 1114 13601 1116
rect 13657 1114 13663 1116
rect 13417 1062 13419 1114
rect 13599 1062 13601 1114
rect 13355 1060 13361 1062
rect 13417 1060 13441 1062
rect 13497 1060 13521 1062
rect 13577 1060 13601 1062
rect 13657 1060 13663 1062
rect 13355 1051 13663 1060
rect 13268 1012 13320 1018
rect 13268 954 13320 960
rect 7656 808 7708 814
rect 7656 750 7708 756
rect 8392 808 8444 814
rect 8392 750 8444 756
rect 10508 808 10560 814
rect 10508 750 10560 756
rect 11428 808 11480 814
rect 11428 750 11480 756
rect 12164 808 12216 814
rect 12164 750 12216 756
rect 13084 808 13136 814
rect 13084 750 13136 756
rect 4100 572 4408 581
rect 4100 570 4106 572
rect 4162 570 4186 572
rect 4242 570 4266 572
rect 4322 570 4346 572
rect 4402 570 4408 572
rect 4162 518 4164 570
rect 4344 518 4346 570
rect 4100 516 4106 518
rect 4162 516 4186 518
rect 4242 516 4266 518
rect 4322 516 4346 518
rect 4402 516 4408 518
rect 4100 507 4408 516
rect 7802 572 8110 581
rect 7802 570 7808 572
rect 7864 570 7888 572
rect 7944 570 7968 572
rect 8024 570 8048 572
rect 8104 570 8110 572
rect 7864 518 7866 570
rect 8046 518 8048 570
rect 7802 516 7808 518
rect 7864 516 7888 518
rect 7944 516 7968 518
rect 8024 516 8048 518
rect 8104 516 8110 518
rect 7802 507 8110 516
rect 8404 474 8432 750
rect 11504 572 11812 581
rect 11504 570 11510 572
rect 11566 570 11590 572
rect 11646 570 11670 572
rect 11726 570 11750 572
rect 11806 570 11812 572
rect 11566 518 11568 570
rect 11748 518 11750 570
rect 11504 516 11510 518
rect 11566 516 11590 518
rect 11646 516 11670 518
rect 11726 516 11750 518
rect 11806 516 11812 518
rect 11504 507 11812 516
rect 15206 572 15514 581
rect 15206 570 15212 572
rect 15268 570 15292 572
rect 15348 570 15372 572
rect 15428 570 15452 572
rect 15508 570 15514 572
rect 15268 518 15270 570
rect 15450 518 15452 570
rect 15206 516 15212 518
rect 15268 516 15292 518
rect 15348 516 15372 518
rect 15428 516 15452 518
rect 15508 516 15514 518
rect 15206 507 15514 516
rect 8024 468 8076 474
rect 7944 428 8024 456
rect 7944 400 7972 428
rect 8024 410 8076 416
rect 8392 468 8444 474
rect 8392 410 8444 416
rect 7930 0 7986 400
<< via2 >>
rect 2255 15258 2311 15260
rect 2335 15258 2391 15260
rect 2415 15258 2471 15260
rect 2495 15258 2551 15260
rect 2255 15206 2301 15258
rect 2301 15206 2311 15258
rect 2335 15206 2365 15258
rect 2365 15206 2377 15258
rect 2377 15206 2391 15258
rect 2415 15206 2429 15258
rect 2429 15206 2441 15258
rect 2441 15206 2471 15258
rect 2495 15206 2505 15258
rect 2505 15206 2551 15258
rect 2255 15204 2311 15206
rect 2335 15204 2391 15206
rect 2415 15204 2471 15206
rect 2495 15204 2551 15206
rect 5957 15258 6013 15260
rect 6037 15258 6093 15260
rect 6117 15258 6173 15260
rect 6197 15258 6253 15260
rect 5957 15206 6003 15258
rect 6003 15206 6013 15258
rect 6037 15206 6067 15258
rect 6067 15206 6079 15258
rect 6079 15206 6093 15258
rect 6117 15206 6131 15258
rect 6131 15206 6143 15258
rect 6143 15206 6173 15258
rect 6197 15206 6207 15258
rect 6207 15206 6253 15258
rect 5957 15204 6013 15206
rect 6037 15204 6093 15206
rect 6117 15204 6173 15206
rect 6197 15204 6253 15206
rect 9659 15258 9715 15260
rect 9739 15258 9795 15260
rect 9819 15258 9875 15260
rect 9899 15258 9955 15260
rect 9659 15206 9705 15258
rect 9705 15206 9715 15258
rect 9739 15206 9769 15258
rect 9769 15206 9781 15258
rect 9781 15206 9795 15258
rect 9819 15206 9833 15258
rect 9833 15206 9845 15258
rect 9845 15206 9875 15258
rect 9899 15206 9909 15258
rect 9909 15206 9955 15258
rect 9659 15204 9715 15206
rect 9739 15204 9795 15206
rect 9819 15204 9875 15206
rect 9899 15204 9955 15206
rect 4106 14714 4162 14716
rect 4186 14714 4242 14716
rect 4266 14714 4322 14716
rect 4346 14714 4402 14716
rect 4106 14662 4152 14714
rect 4152 14662 4162 14714
rect 4186 14662 4216 14714
rect 4216 14662 4228 14714
rect 4228 14662 4242 14714
rect 4266 14662 4280 14714
rect 4280 14662 4292 14714
rect 4292 14662 4322 14714
rect 4346 14662 4356 14714
rect 4356 14662 4402 14714
rect 4106 14660 4162 14662
rect 4186 14660 4242 14662
rect 4266 14660 4322 14662
rect 4346 14660 4402 14662
rect 7808 14714 7864 14716
rect 7888 14714 7944 14716
rect 7968 14714 8024 14716
rect 8048 14714 8104 14716
rect 7808 14662 7854 14714
rect 7854 14662 7864 14714
rect 7888 14662 7918 14714
rect 7918 14662 7930 14714
rect 7930 14662 7944 14714
rect 7968 14662 7982 14714
rect 7982 14662 7994 14714
rect 7994 14662 8024 14714
rect 8048 14662 8058 14714
rect 8058 14662 8104 14714
rect 7808 14660 7864 14662
rect 7888 14660 7944 14662
rect 7968 14660 8024 14662
rect 8048 14660 8104 14662
rect 2255 14170 2311 14172
rect 2335 14170 2391 14172
rect 2415 14170 2471 14172
rect 2495 14170 2551 14172
rect 2255 14118 2301 14170
rect 2301 14118 2311 14170
rect 2335 14118 2365 14170
rect 2365 14118 2377 14170
rect 2377 14118 2391 14170
rect 2415 14118 2429 14170
rect 2429 14118 2441 14170
rect 2441 14118 2471 14170
rect 2495 14118 2505 14170
rect 2505 14118 2551 14170
rect 2255 14116 2311 14118
rect 2335 14116 2391 14118
rect 2415 14116 2471 14118
rect 2495 14116 2551 14118
rect 5957 14170 6013 14172
rect 6037 14170 6093 14172
rect 6117 14170 6173 14172
rect 6197 14170 6253 14172
rect 5957 14118 6003 14170
rect 6003 14118 6013 14170
rect 6037 14118 6067 14170
rect 6067 14118 6079 14170
rect 6079 14118 6093 14170
rect 6117 14118 6131 14170
rect 6131 14118 6143 14170
rect 6143 14118 6173 14170
rect 6197 14118 6207 14170
rect 6207 14118 6253 14170
rect 5957 14116 6013 14118
rect 6037 14116 6093 14118
rect 6117 14116 6173 14118
rect 6197 14116 6253 14118
rect 11510 14714 11566 14716
rect 11590 14714 11646 14716
rect 11670 14714 11726 14716
rect 11750 14714 11806 14716
rect 11510 14662 11556 14714
rect 11556 14662 11566 14714
rect 11590 14662 11620 14714
rect 11620 14662 11632 14714
rect 11632 14662 11646 14714
rect 11670 14662 11684 14714
rect 11684 14662 11696 14714
rect 11696 14662 11726 14714
rect 11750 14662 11760 14714
rect 11760 14662 11806 14714
rect 11510 14660 11566 14662
rect 11590 14660 11646 14662
rect 11670 14660 11726 14662
rect 11750 14660 11806 14662
rect 9659 14170 9715 14172
rect 9739 14170 9795 14172
rect 9819 14170 9875 14172
rect 9899 14170 9955 14172
rect 9659 14118 9705 14170
rect 9705 14118 9715 14170
rect 9739 14118 9769 14170
rect 9769 14118 9781 14170
rect 9781 14118 9795 14170
rect 9819 14118 9833 14170
rect 9833 14118 9845 14170
rect 9845 14118 9875 14170
rect 9899 14118 9909 14170
rect 9909 14118 9955 14170
rect 9659 14116 9715 14118
rect 9739 14116 9795 14118
rect 9819 14116 9875 14118
rect 9899 14116 9955 14118
rect 4106 13626 4162 13628
rect 4186 13626 4242 13628
rect 4266 13626 4322 13628
rect 4346 13626 4402 13628
rect 4106 13574 4152 13626
rect 4152 13574 4162 13626
rect 4186 13574 4216 13626
rect 4216 13574 4228 13626
rect 4228 13574 4242 13626
rect 4266 13574 4280 13626
rect 4280 13574 4292 13626
rect 4292 13574 4322 13626
rect 4346 13574 4356 13626
rect 4356 13574 4402 13626
rect 4106 13572 4162 13574
rect 4186 13572 4242 13574
rect 4266 13572 4322 13574
rect 4346 13572 4402 13574
rect 7808 13626 7864 13628
rect 7888 13626 7944 13628
rect 7968 13626 8024 13628
rect 8048 13626 8104 13628
rect 7808 13574 7854 13626
rect 7854 13574 7864 13626
rect 7888 13574 7918 13626
rect 7918 13574 7930 13626
rect 7930 13574 7944 13626
rect 7968 13574 7982 13626
rect 7982 13574 7994 13626
rect 7994 13574 8024 13626
rect 8048 13574 8058 13626
rect 8058 13574 8104 13626
rect 7808 13572 7864 13574
rect 7888 13572 7944 13574
rect 7968 13572 8024 13574
rect 8048 13572 8104 13574
rect 11510 13626 11566 13628
rect 11590 13626 11646 13628
rect 11670 13626 11726 13628
rect 11750 13626 11806 13628
rect 11510 13574 11556 13626
rect 11556 13574 11566 13626
rect 11590 13574 11620 13626
rect 11620 13574 11632 13626
rect 11632 13574 11646 13626
rect 11670 13574 11684 13626
rect 11684 13574 11696 13626
rect 11696 13574 11726 13626
rect 11750 13574 11760 13626
rect 11760 13574 11806 13626
rect 11510 13572 11566 13574
rect 11590 13572 11646 13574
rect 11670 13572 11726 13574
rect 11750 13572 11806 13574
rect 2255 13082 2311 13084
rect 2335 13082 2391 13084
rect 2415 13082 2471 13084
rect 2495 13082 2551 13084
rect 2255 13030 2301 13082
rect 2301 13030 2311 13082
rect 2335 13030 2365 13082
rect 2365 13030 2377 13082
rect 2377 13030 2391 13082
rect 2415 13030 2429 13082
rect 2429 13030 2441 13082
rect 2441 13030 2471 13082
rect 2495 13030 2505 13082
rect 2505 13030 2551 13082
rect 2255 13028 2311 13030
rect 2335 13028 2391 13030
rect 2415 13028 2471 13030
rect 2495 13028 2551 13030
rect 5957 13082 6013 13084
rect 6037 13082 6093 13084
rect 6117 13082 6173 13084
rect 6197 13082 6253 13084
rect 5957 13030 6003 13082
rect 6003 13030 6013 13082
rect 6037 13030 6067 13082
rect 6067 13030 6079 13082
rect 6079 13030 6093 13082
rect 6117 13030 6131 13082
rect 6131 13030 6143 13082
rect 6143 13030 6173 13082
rect 6197 13030 6207 13082
rect 6207 13030 6253 13082
rect 5957 13028 6013 13030
rect 6037 13028 6093 13030
rect 6117 13028 6173 13030
rect 6197 13028 6253 13030
rect 4106 12538 4162 12540
rect 4186 12538 4242 12540
rect 4266 12538 4322 12540
rect 4346 12538 4402 12540
rect 4106 12486 4152 12538
rect 4152 12486 4162 12538
rect 4186 12486 4216 12538
rect 4216 12486 4228 12538
rect 4228 12486 4242 12538
rect 4266 12486 4280 12538
rect 4280 12486 4292 12538
rect 4292 12486 4322 12538
rect 4346 12486 4356 12538
rect 4356 12486 4402 12538
rect 4106 12484 4162 12486
rect 4186 12484 4242 12486
rect 4266 12484 4322 12486
rect 4346 12484 4402 12486
rect 7808 12538 7864 12540
rect 7888 12538 7944 12540
rect 7968 12538 8024 12540
rect 8048 12538 8104 12540
rect 7808 12486 7854 12538
rect 7854 12486 7864 12538
rect 7888 12486 7918 12538
rect 7918 12486 7930 12538
rect 7930 12486 7944 12538
rect 7968 12486 7982 12538
rect 7982 12486 7994 12538
rect 7994 12486 8024 12538
rect 8048 12486 8058 12538
rect 8058 12486 8104 12538
rect 7808 12484 7864 12486
rect 7888 12484 7944 12486
rect 7968 12484 8024 12486
rect 8048 12484 8104 12486
rect 9659 13082 9715 13084
rect 9739 13082 9795 13084
rect 9819 13082 9875 13084
rect 9899 13082 9955 13084
rect 9659 13030 9705 13082
rect 9705 13030 9715 13082
rect 9739 13030 9769 13082
rect 9769 13030 9781 13082
rect 9781 13030 9795 13082
rect 9819 13030 9833 13082
rect 9833 13030 9845 13082
rect 9845 13030 9875 13082
rect 9899 13030 9909 13082
rect 9909 13030 9955 13082
rect 9659 13028 9715 13030
rect 9739 13028 9795 13030
rect 9819 13028 9875 13030
rect 9899 13028 9955 13030
rect 2255 11994 2311 11996
rect 2335 11994 2391 11996
rect 2415 11994 2471 11996
rect 2495 11994 2551 11996
rect 2255 11942 2301 11994
rect 2301 11942 2311 11994
rect 2335 11942 2365 11994
rect 2365 11942 2377 11994
rect 2377 11942 2391 11994
rect 2415 11942 2429 11994
rect 2429 11942 2441 11994
rect 2441 11942 2471 11994
rect 2495 11942 2505 11994
rect 2505 11942 2551 11994
rect 2255 11940 2311 11942
rect 2335 11940 2391 11942
rect 2415 11940 2471 11942
rect 2495 11940 2551 11942
rect 5957 11994 6013 11996
rect 6037 11994 6093 11996
rect 6117 11994 6173 11996
rect 6197 11994 6253 11996
rect 5957 11942 6003 11994
rect 6003 11942 6013 11994
rect 6037 11942 6067 11994
rect 6067 11942 6079 11994
rect 6079 11942 6093 11994
rect 6117 11942 6131 11994
rect 6131 11942 6143 11994
rect 6143 11942 6173 11994
rect 6197 11942 6207 11994
rect 6207 11942 6253 11994
rect 5957 11940 6013 11942
rect 6037 11940 6093 11942
rect 6117 11940 6173 11942
rect 6197 11940 6253 11942
rect 4106 11450 4162 11452
rect 4186 11450 4242 11452
rect 4266 11450 4322 11452
rect 4346 11450 4402 11452
rect 4106 11398 4152 11450
rect 4152 11398 4162 11450
rect 4186 11398 4216 11450
rect 4216 11398 4228 11450
rect 4228 11398 4242 11450
rect 4266 11398 4280 11450
rect 4280 11398 4292 11450
rect 4292 11398 4322 11450
rect 4346 11398 4356 11450
rect 4356 11398 4402 11450
rect 4106 11396 4162 11398
rect 4186 11396 4242 11398
rect 4266 11396 4322 11398
rect 4346 11396 4402 11398
rect 7808 11450 7864 11452
rect 7888 11450 7944 11452
rect 7968 11450 8024 11452
rect 8048 11450 8104 11452
rect 7808 11398 7854 11450
rect 7854 11398 7864 11450
rect 7888 11398 7918 11450
rect 7918 11398 7930 11450
rect 7930 11398 7944 11450
rect 7968 11398 7982 11450
rect 7982 11398 7994 11450
rect 7994 11398 8024 11450
rect 8048 11398 8058 11450
rect 8058 11398 8104 11450
rect 7808 11396 7864 11398
rect 7888 11396 7944 11398
rect 7968 11396 8024 11398
rect 8048 11396 8104 11398
rect 2255 10906 2311 10908
rect 2335 10906 2391 10908
rect 2415 10906 2471 10908
rect 2495 10906 2551 10908
rect 2255 10854 2301 10906
rect 2301 10854 2311 10906
rect 2335 10854 2365 10906
rect 2365 10854 2377 10906
rect 2377 10854 2391 10906
rect 2415 10854 2429 10906
rect 2429 10854 2441 10906
rect 2441 10854 2471 10906
rect 2495 10854 2505 10906
rect 2505 10854 2551 10906
rect 2255 10852 2311 10854
rect 2335 10852 2391 10854
rect 2415 10852 2471 10854
rect 2495 10852 2551 10854
rect 5957 10906 6013 10908
rect 6037 10906 6093 10908
rect 6117 10906 6173 10908
rect 6197 10906 6253 10908
rect 5957 10854 6003 10906
rect 6003 10854 6013 10906
rect 6037 10854 6067 10906
rect 6067 10854 6079 10906
rect 6079 10854 6093 10906
rect 6117 10854 6131 10906
rect 6131 10854 6143 10906
rect 6143 10854 6173 10906
rect 6197 10854 6207 10906
rect 6207 10854 6253 10906
rect 5957 10852 6013 10854
rect 6037 10852 6093 10854
rect 6117 10852 6173 10854
rect 6197 10852 6253 10854
rect 4106 10362 4162 10364
rect 4186 10362 4242 10364
rect 4266 10362 4322 10364
rect 4346 10362 4402 10364
rect 4106 10310 4152 10362
rect 4152 10310 4162 10362
rect 4186 10310 4216 10362
rect 4216 10310 4228 10362
rect 4228 10310 4242 10362
rect 4266 10310 4280 10362
rect 4280 10310 4292 10362
rect 4292 10310 4322 10362
rect 4346 10310 4356 10362
rect 4356 10310 4402 10362
rect 4106 10308 4162 10310
rect 4186 10308 4242 10310
rect 4266 10308 4322 10310
rect 4346 10308 4402 10310
rect 7808 10362 7864 10364
rect 7888 10362 7944 10364
rect 7968 10362 8024 10364
rect 8048 10362 8104 10364
rect 7808 10310 7854 10362
rect 7854 10310 7864 10362
rect 7888 10310 7918 10362
rect 7918 10310 7930 10362
rect 7930 10310 7944 10362
rect 7968 10310 7982 10362
rect 7982 10310 7994 10362
rect 7994 10310 8024 10362
rect 8048 10310 8058 10362
rect 8058 10310 8104 10362
rect 7808 10308 7864 10310
rect 7888 10308 7944 10310
rect 7968 10308 8024 10310
rect 8048 10308 8104 10310
rect 2255 9818 2311 9820
rect 2335 9818 2391 9820
rect 2415 9818 2471 9820
rect 2495 9818 2551 9820
rect 2255 9766 2301 9818
rect 2301 9766 2311 9818
rect 2335 9766 2365 9818
rect 2365 9766 2377 9818
rect 2377 9766 2391 9818
rect 2415 9766 2429 9818
rect 2429 9766 2441 9818
rect 2441 9766 2471 9818
rect 2495 9766 2505 9818
rect 2505 9766 2551 9818
rect 2255 9764 2311 9766
rect 2335 9764 2391 9766
rect 2415 9764 2471 9766
rect 2495 9764 2551 9766
rect 5957 9818 6013 9820
rect 6037 9818 6093 9820
rect 6117 9818 6173 9820
rect 6197 9818 6253 9820
rect 5957 9766 6003 9818
rect 6003 9766 6013 9818
rect 6037 9766 6067 9818
rect 6067 9766 6079 9818
rect 6079 9766 6093 9818
rect 6117 9766 6131 9818
rect 6131 9766 6143 9818
rect 6143 9766 6173 9818
rect 6197 9766 6207 9818
rect 6207 9766 6253 9818
rect 5957 9764 6013 9766
rect 6037 9764 6093 9766
rect 6117 9764 6173 9766
rect 6197 9764 6253 9766
rect 4106 9274 4162 9276
rect 4186 9274 4242 9276
rect 4266 9274 4322 9276
rect 4346 9274 4402 9276
rect 4106 9222 4152 9274
rect 4152 9222 4162 9274
rect 4186 9222 4216 9274
rect 4216 9222 4228 9274
rect 4228 9222 4242 9274
rect 4266 9222 4280 9274
rect 4280 9222 4292 9274
rect 4292 9222 4322 9274
rect 4346 9222 4356 9274
rect 4356 9222 4402 9274
rect 4106 9220 4162 9222
rect 4186 9220 4242 9222
rect 4266 9220 4322 9222
rect 4346 9220 4402 9222
rect 7808 9274 7864 9276
rect 7888 9274 7944 9276
rect 7968 9274 8024 9276
rect 8048 9274 8104 9276
rect 7808 9222 7854 9274
rect 7854 9222 7864 9274
rect 7888 9222 7918 9274
rect 7918 9222 7930 9274
rect 7930 9222 7944 9274
rect 7968 9222 7982 9274
rect 7982 9222 7994 9274
rect 7994 9222 8024 9274
rect 8048 9222 8058 9274
rect 8058 9222 8104 9274
rect 7808 9220 7864 9222
rect 7888 9220 7944 9222
rect 7968 9220 8024 9222
rect 8048 9220 8104 9222
rect 9659 11994 9715 11996
rect 9739 11994 9795 11996
rect 9819 11994 9875 11996
rect 9899 11994 9955 11996
rect 9659 11942 9705 11994
rect 9705 11942 9715 11994
rect 9739 11942 9769 11994
rect 9769 11942 9781 11994
rect 9781 11942 9795 11994
rect 9819 11942 9833 11994
rect 9833 11942 9845 11994
rect 9845 11942 9875 11994
rect 9899 11942 9909 11994
rect 9909 11942 9955 11994
rect 9659 11940 9715 11942
rect 9739 11940 9795 11942
rect 9819 11940 9875 11942
rect 9899 11940 9955 11942
rect 11510 12538 11566 12540
rect 11590 12538 11646 12540
rect 11670 12538 11726 12540
rect 11750 12538 11806 12540
rect 11510 12486 11556 12538
rect 11556 12486 11566 12538
rect 11590 12486 11620 12538
rect 11620 12486 11632 12538
rect 11632 12486 11646 12538
rect 11670 12486 11684 12538
rect 11684 12486 11696 12538
rect 11696 12486 11726 12538
rect 11750 12486 11760 12538
rect 11760 12486 11806 12538
rect 11510 12484 11566 12486
rect 11590 12484 11646 12486
rect 11670 12484 11726 12486
rect 11750 12484 11806 12486
rect 11510 11450 11566 11452
rect 11590 11450 11646 11452
rect 11670 11450 11726 11452
rect 11750 11450 11806 11452
rect 11510 11398 11556 11450
rect 11556 11398 11566 11450
rect 11590 11398 11620 11450
rect 11620 11398 11632 11450
rect 11632 11398 11646 11450
rect 11670 11398 11684 11450
rect 11684 11398 11696 11450
rect 11696 11398 11726 11450
rect 11750 11398 11760 11450
rect 11760 11398 11806 11450
rect 11510 11396 11566 11398
rect 11590 11396 11646 11398
rect 11670 11396 11726 11398
rect 11750 11396 11806 11398
rect 2255 8730 2311 8732
rect 2335 8730 2391 8732
rect 2415 8730 2471 8732
rect 2495 8730 2551 8732
rect 2255 8678 2301 8730
rect 2301 8678 2311 8730
rect 2335 8678 2365 8730
rect 2365 8678 2377 8730
rect 2377 8678 2391 8730
rect 2415 8678 2429 8730
rect 2429 8678 2441 8730
rect 2441 8678 2471 8730
rect 2495 8678 2505 8730
rect 2505 8678 2551 8730
rect 2255 8676 2311 8678
rect 2335 8676 2391 8678
rect 2415 8676 2471 8678
rect 2495 8676 2551 8678
rect 5957 8730 6013 8732
rect 6037 8730 6093 8732
rect 6117 8730 6173 8732
rect 6197 8730 6253 8732
rect 5957 8678 6003 8730
rect 6003 8678 6013 8730
rect 6037 8678 6067 8730
rect 6067 8678 6079 8730
rect 6079 8678 6093 8730
rect 6117 8678 6131 8730
rect 6131 8678 6143 8730
rect 6143 8678 6173 8730
rect 6197 8678 6207 8730
rect 6207 8678 6253 8730
rect 5957 8676 6013 8678
rect 6037 8676 6093 8678
rect 6117 8676 6173 8678
rect 6197 8676 6253 8678
rect 4106 8186 4162 8188
rect 4186 8186 4242 8188
rect 4266 8186 4322 8188
rect 4346 8186 4402 8188
rect 4106 8134 4152 8186
rect 4152 8134 4162 8186
rect 4186 8134 4216 8186
rect 4216 8134 4228 8186
rect 4228 8134 4242 8186
rect 4266 8134 4280 8186
rect 4280 8134 4292 8186
rect 4292 8134 4322 8186
rect 4346 8134 4356 8186
rect 4356 8134 4402 8186
rect 4106 8132 4162 8134
rect 4186 8132 4242 8134
rect 4266 8132 4322 8134
rect 4346 8132 4402 8134
rect 7808 8186 7864 8188
rect 7888 8186 7944 8188
rect 7968 8186 8024 8188
rect 8048 8186 8104 8188
rect 7808 8134 7854 8186
rect 7854 8134 7864 8186
rect 7888 8134 7918 8186
rect 7918 8134 7930 8186
rect 7930 8134 7944 8186
rect 7968 8134 7982 8186
rect 7982 8134 7994 8186
rect 7994 8134 8024 8186
rect 8048 8134 8058 8186
rect 8058 8134 8104 8186
rect 7808 8132 7864 8134
rect 7888 8132 7944 8134
rect 7968 8132 8024 8134
rect 8048 8132 8104 8134
rect 9659 10906 9715 10908
rect 9739 10906 9795 10908
rect 9819 10906 9875 10908
rect 9899 10906 9955 10908
rect 9659 10854 9705 10906
rect 9705 10854 9715 10906
rect 9739 10854 9769 10906
rect 9769 10854 9781 10906
rect 9781 10854 9795 10906
rect 9819 10854 9833 10906
rect 9833 10854 9845 10906
rect 9845 10854 9875 10906
rect 9899 10854 9909 10906
rect 9909 10854 9955 10906
rect 9659 10852 9715 10854
rect 9739 10852 9795 10854
rect 9819 10852 9875 10854
rect 9899 10852 9955 10854
rect 9659 9818 9715 9820
rect 9739 9818 9795 9820
rect 9819 9818 9875 9820
rect 9899 9818 9955 9820
rect 9659 9766 9705 9818
rect 9705 9766 9715 9818
rect 9739 9766 9769 9818
rect 9769 9766 9781 9818
rect 9781 9766 9795 9818
rect 9819 9766 9833 9818
rect 9833 9766 9845 9818
rect 9845 9766 9875 9818
rect 9899 9766 9909 9818
rect 9909 9766 9955 9818
rect 9659 9764 9715 9766
rect 9739 9764 9795 9766
rect 9819 9764 9875 9766
rect 9899 9764 9955 9766
rect 9218 7964 9220 7984
rect 9220 7964 9272 7984
rect 9272 7964 9274 7984
rect 9218 7928 9274 7964
rect 2255 7642 2311 7644
rect 2335 7642 2391 7644
rect 2415 7642 2471 7644
rect 2495 7642 2551 7644
rect 2255 7590 2301 7642
rect 2301 7590 2311 7642
rect 2335 7590 2365 7642
rect 2365 7590 2377 7642
rect 2377 7590 2391 7642
rect 2415 7590 2429 7642
rect 2429 7590 2441 7642
rect 2441 7590 2471 7642
rect 2495 7590 2505 7642
rect 2505 7590 2551 7642
rect 2255 7588 2311 7590
rect 2335 7588 2391 7590
rect 2415 7588 2471 7590
rect 2495 7588 2551 7590
rect 5957 7642 6013 7644
rect 6037 7642 6093 7644
rect 6117 7642 6173 7644
rect 6197 7642 6253 7644
rect 5957 7590 6003 7642
rect 6003 7590 6013 7642
rect 6037 7590 6067 7642
rect 6067 7590 6079 7642
rect 6079 7590 6093 7642
rect 6117 7590 6131 7642
rect 6131 7590 6143 7642
rect 6143 7590 6173 7642
rect 6197 7590 6207 7642
rect 6207 7590 6253 7642
rect 5957 7588 6013 7590
rect 6037 7588 6093 7590
rect 6117 7588 6173 7590
rect 6197 7588 6253 7590
rect 4106 7098 4162 7100
rect 4186 7098 4242 7100
rect 4266 7098 4322 7100
rect 4346 7098 4402 7100
rect 4106 7046 4152 7098
rect 4152 7046 4162 7098
rect 4186 7046 4216 7098
rect 4216 7046 4228 7098
rect 4228 7046 4242 7098
rect 4266 7046 4280 7098
rect 4280 7046 4292 7098
rect 4292 7046 4322 7098
rect 4346 7046 4356 7098
rect 4356 7046 4402 7098
rect 4106 7044 4162 7046
rect 4186 7044 4242 7046
rect 4266 7044 4322 7046
rect 4346 7044 4402 7046
rect 7808 7098 7864 7100
rect 7888 7098 7944 7100
rect 7968 7098 8024 7100
rect 8048 7098 8104 7100
rect 7808 7046 7854 7098
rect 7854 7046 7864 7098
rect 7888 7046 7918 7098
rect 7918 7046 7930 7098
rect 7930 7046 7944 7098
rect 7968 7046 7982 7098
rect 7982 7046 7994 7098
rect 7994 7046 8024 7098
rect 8048 7046 8058 7098
rect 8058 7046 8104 7098
rect 7808 7044 7864 7046
rect 7888 7044 7944 7046
rect 7968 7044 8024 7046
rect 8048 7044 8104 7046
rect 2255 6554 2311 6556
rect 2335 6554 2391 6556
rect 2415 6554 2471 6556
rect 2495 6554 2551 6556
rect 2255 6502 2301 6554
rect 2301 6502 2311 6554
rect 2335 6502 2365 6554
rect 2365 6502 2377 6554
rect 2377 6502 2391 6554
rect 2415 6502 2429 6554
rect 2429 6502 2441 6554
rect 2441 6502 2471 6554
rect 2495 6502 2505 6554
rect 2505 6502 2551 6554
rect 2255 6500 2311 6502
rect 2335 6500 2391 6502
rect 2415 6500 2471 6502
rect 2495 6500 2551 6502
rect 5957 6554 6013 6556
rect 6037 6554 6093 6556
rect 6117 6554 6173 6556
rect 6197 6554 6253 6556
rect 5957 6502 6003 6554
rect 6003 6502 6013 6554
rect 6037 6502 6067 6554
rect 6067 6502 6079 6554
rect 6079 6502 6093 6554
rect 6117 6502 6131 6554
rect 6131 6502 6143 6554
rect 6143 6502 6173 6554
rect 6197 6502 6207 6554
rect 6207 6502 6253 6554
rect 5957 6500 6013 6502
rect 6037 6500 6093 6502
rect 6117 6500 6173 6502
rect 6197 6500 6253 6502
rect 4106 6010 4162 6012
rect 4186 6010 4242 6012
rect 4266 6010 4322 6012
rect 4346 6010 4402 6012
rect 4106 5958 4152 6010
rect 4152 5958 4162 6010
rect 4186 5958 4216 6010
rect 4216 5958 4228 6010
rect 4228 5958 4242 6010
rect 4266 5958 4280 6010
rect 4280 5958 4292 6010
rect 4292 5958 4322 6010
rect 4346 5958 4356 6010
rect 4356 5958 4402 6010
rect 4106 5956 4162 5958
rect 4186 5956 4242 5958
rect 4266 5956 4322 5958
rect 4346 5956 4402 5958
rect 7808 6010 7864 6012
rect 7888 6010 7944 6012
rect 7968 6010 8024 6012
rect 8048 6010 8104 6012
rect 7808 5958 7854 6010
rect 7854 5958 7864 6010
rect 7888 5958 7918 6010
rect 7918 5958 7930 6010
rect 7930 5958 7944 6010
rect 7968 5958 7982 6010
rect 7982 5958 7994 6010
rect 7994 5958 8024 6010
rect 8048 5958 8058 6010
rect 8058 5958 8104 6010
rect 7808 5956 7864 5958
rect 7888 5956 7944 5958
rect 7968 5956 8024 5958
rect 8048 5956 8104 5958
rect 2255 5466 2311 5468
rect 2335 5466 2391 5468
rect 2415 5466 2471 5468
rect 2495 5466 2551 5468
rect 2255 5414 2301 5466
rect 2301 5414 2311 5466
rect 2335 5414 2365 5466
rect 2365 5414 2377 5466
rect 2377 5414 2391 5466
rect 2415 5414 2429 5466
rect 2429 5414 2441 5466
rect 2441 5414 2471 5466
rect 2495 5414 2505 5466
rect 2505 5414 2551 5466
rect 2255 5412 2311 5414
rect 2335 5412 2391 5414
rect 2415 5412 2471 5414
rect 2495 5412 2551 5414
rect 5957 5466 6013 5468
rect 6037 5466 6093 5468
rect 6117 5466 6173 5468
rect 6197 5466 6253 5468
rect 5957 5414 6003 5466
rect 6003 5414 6013 5466
rect 6037 5414 6067 5466
rect 6067 5414 6079 5466
rect 6079 5414 6093 5466
rect 6117 5414 6131 5466
rect 6131 5414 6143 5466
rect 6143 5414 6173 5466
rect 6197 5414 6207 5466
rect 6207 5414 6253 5466
rect 5957 5412 6013 5414
rect 6037 5412 6093 5414
rect 6117 5412 6173 5414
rect 6197 5412 6253 5414
rect 8390 5752 8446 5808
rect 9770 9036 9826 9072
rect 9770 9016 9772 9036
rect 9772 9016 9824 9036
rect 9824 9016 9826 9036
rect 10506 9036 10562 9072
rect 10506 9016 10508 9036
rect 10508 9016 10560 9036
rect 10560 9016 10562 9036
rect 9659 8730 9715 8732
rect 9739 8730 9795 8732
rect 9819 8730 9875 8732
rect 9899 8730 9955 8732
rect 9659 8678 9705 8730
rect 9705 8678 9715 8730
rect 9739 8678 9769 8730
rect 9769 8678 9781 8730
rect 9781 8678 9795 8730
rect 9819 8678 9833 8730
rect 9833 8678 9845 8730
rect 9845 8678 9875 8730
rect 9899 8678 9909 8730
rect 9909 8678 9955 8730
rect 9659 8676 9715 8678
rect 9739 8676 9795 8678
rect 9819 8676 9875 8678
rect 9899 8676 9955 8678
rect 11510 10362 11566 10364
rect 11590 10362 11646 10364
rect 11670 10362 11726 10364
rect 11750 10362 11806 10364
rect 11510 10310 11556 10362
rect 11556 10310 11566 10362
rect 11590 10310 11620 10362
rect 11620 10310 11632 10362
rect 11632 10310 11646 10362
rect 11670 10310 11684 10362
rect 11684 10310 11696 10362
rect 11696 10310 11726 10362
rect 11750 10310 11760 10362
rect 11760 10310 11806 10362
rect 11510 10308 11566 10310
rect 11590 10308 11646 10310
rect 11670 10308 11726 10310
rect 11750 10308 11806 10310
rect 11510 9274 11566 9276
rect 11590 9274 11646 9276
rect 11670 9274 11726 9276
rect 11750 9274 11806 9276
rect 11510 9222 11556 9274
rect 11556 9222 11566 9274
rect 11590 9222 11620 9274
rect 11620 9222 11632 9274
rect 11632 9222 11646 9274
rect 11670 9222 11684 9274
rect 11684 9222 11696 9274
rect 11696 9222 11726 9274
rect 11750 9222 11760 9274
rect 11760 9222 11806 9274
rect 11510 9220 11566 9222
rect 11590 9220 11646 9222
rect 11670 9220 11726 9222
rect 11750 9220 11806 9222
rect 9659 7642 9715 7644
rect 9739 7642 9795 7644
rect 9819 7642 9875 7644
rect 9899 7642 9955 7644
rect 9659 7590 9705 7642
rect 9705 7590 9715 7642
rect 9739 7590 9769 7642
rect 9769 7590 9781 7642
rect 9781 7590 9795 7642
rect 9819 7590 9833 7642
rect 9833 7590 9845 7642
rect 9845 7590 9875 7642
rect 9899 7590 9909 7642
rect 9909 7590 9955 7642
rect 9659 7588 9715 7590
rect 9739 7588 9795 7590
rect 9819 7588 9875 7590
rect 9899 7588 9955 7590
rect 9218 6840 9274 6896
rect 4106 4922 4162 4924
rect 4186 4922 4242 4924
rect 4266 4922 4322 4924
rect 4346 4922 4402 4924
rect 4106 4870 4152 4922
rect 4152 4870 4162 4922
rect 4186 4870 4216 4922
rect 4216 4870 4228 4922
rect 4228 4870 4242 4922
rect 4266 4870 4280 4922
rect 4280 4870 4292 4922
rect 4292 4870 4322 4922
rect 4346 4870 4356 4922
rect 4356 4870 4402 4922
rect 4106 4868 4162 4870
rect 4186 4868 4242 4870
rect 4266 4868 4322 4870
rect 4346 4868 4402 4870
rect 7808 4922 7864 4924
rect 7888 4922 7944 4924
rect 7968 4922 8024 4924
rect 8048 4922 8104 4924
rect 7808 4870 7854 4922
rect 7854 4870 7864 4922
rect 7888 4870 7918 4922
rect 7918 4870 7930 4922
rect 7930 4870 7944 4922
rect 7968 4870 7982 4922
rect 7982 4870 7994 4922
rect 7994 4870 8024 4922
rect 8048 4870 8058 4922
rect 8058 4870 8104 4922
rect 7808 4868 7864 4870
rect 7888 4868 7944 4870
rect 7968 4868 8024 4870
rect 8048 4868 8104 4870
rect 2255 4378 2311 4380
rect 2335 4378 2391 4380
rect 2415 4378 2471 4380
rect 2495 4378 2551 4380
rect 2255 4326 2301 4378
rect 2301 4326 2311 4378
rect 2335 4326 2365 4378
rect 2365 4326 2377 4378
rect 2377 4326 2391 4378
rect 2415 4326 2429 4378
rect 2429 4326 2441 4378
rect 2441 4326 2471 4378
rect 2495 4326 2505 4378
rect 2505 4326 2551 4378
rect 2255 4324 2311 4326
rect 2335 4324 2391 4326
rect 2415 4324 2471 4326
rect 2495 4324 2551 4326
rect 5957 4378 6013 4380
rect 6037 4378 6093 4380
rect 6117 4378 6173 4380
rect 6197 4378 6253 4380
rect 5957 4326 6003 4378
rect 6003 4326 6013 4378
rect 6037 4326 6067 4378
rect 6067 4326 6079 4378
rect 6079 4326 6093 4378
rect 6117 4326 6131 4378
rect 6131 4326 6143 4378
rect 6143 4326 6173 4378
rect 6197 4326 6207 4378
rect 6207 4326 6253 4378
rect 5957 4324 6013 4326
rect 6037 4324 6093 4326
rect 6117 4324 6173 4326
rect 6197 4324 6253 4326
rect 4106 3834 4162 3836
rect 4186 3834 4242 3836
rect 4266 3834 4322 3836
rect 4346 3834 4402 3836
rect 4106 3782 4152 3834
rect 4152 3782 4162 3834
rect 4186 3782 4216 3834
rect 4216 3782 4228 3834
rect 4228 3782 4242 3834
rect 4266 3782 4280 3834
rect 4280 3782 4292 3834
rect 4292 3782 4322 3834
rect 4346 3782 4356 3834
rect 4356 3782 4402 3834
rect 4106 3780 4162 3782
rect 4186 3780 4242 3782
rect 4266 3780 4322 3782
rect 4346 3780 4402 3782
rect 2255 3290 2311 3292
rect 2335 3290 2391 3292
rect 2415 3290 2471 3292
rect 2495 3290 2551 3292
rect 2255 3238 2301 3290
rect 2301 3238 2311 3290
rect 2335 3238 2365 3290
rect 2365 3238 2377 3290
rect 2377 3238 2391 3290
rect 2415 3238 2429 3290
rect 2429 3238 2441 3290
rect 2441 3238 2471 3290
rect 2495 3238 2505 3290
rect 2505 3238 2551 3290
rect 2255 3236 2311 3238
rect 2335 3236 2391 3238
rect 2415 3236 2471 3238
rect 2495 3236 2551 3238
rect 5957 3290 6013 3292
rect 6037 3290 6093 3292
rect 6117 3290 6173 3292
rect 6197 3290 6253 3292
rect 5957 3238 6003 3290
rect 6003 3238 6013 3290
rect 6037 3238 6067 3290
rect 6067 3238 6079 3290
rect 6079 3238 6093 3290
rect 6117 3238 6131 3290
rect 6131 3238 6143 3290
rect 6143 3238 6173 3290
rect 6197 3238 6207 3290
rect 6207 3238 6253 3290
rect 5957 3236 6013 3238
rect 6037 3236 6093 3238
rect 6117 3236 6173 3238
rect 6197 3236 6253 3238
rect 7808 3834 7864 3836
rect 7888 3834 7944 3836
rect 7968 3834 8024 3836
rect 8048 3834 8104 3836
rect 7808 3782 7854 3834
rect 7854 3782 7864 3834
rect 7888 3782 7918 3834
rect 7918 3782 7930 3834
rect 7930 3782 7944 3834
rect 7968 3782 7982 3834
rect 7982 3782 7994 3834
rect 7994 3782 8024 3834
rect 8048 3782 8058 3834
rect 8058 3782 8104 3834
rect 7808 3780 7864 3782
rect 7888 3780 7944 3782
rect 7968 3780 8024 3782
rect 8048 3780 8104 3782
rect 9659 6554 9715 6556
rect 9739 6554 9795 6556
rect 9819 6554 9875 6556
rect 9899 6554 9955 6556
rect 9659 6502 9705 6554
rect 9705 6502 9715 6554
rect 9739 6502 9769 6554
rect 9769 6502 9781 6554
rect 9781 6502 9795 6554
rect 9819 6502 9833 6554
rect 9833 6502 9845 6554
rect 9845 6502 9875 6554
rect 9899 6502 9909 6554
rect 9909 6502 9955 6554
rect 9659 6500 9715 6502
rect 9739 6500 9795 6502
rect 9819 6500 9875 6502
rect 9899 6500 9955 6502
rect 11510 8186 11566 8188
rect 11590 8186 11646 8188
rect 11670 8186 11726 8188
rect 11750 8186 11806 8188
rect 11510 8134 11556 8186
rect 11556 8134 11566 8186
rect 11590 8134 11620 8186
rect 11620 8134 11632 8186
rect 11632 8134 11646 8186
rect 11670 8134 11684 8186
rect 11684 8134 11696 8186
rect 11696 8134 11726 8186
rect 11750 8134 11760 8186
rect 11760 8134 11806 8186
rect 11510 8132 11566 8134
rect 11590 8132 11646 8134
rect 11670 8132 11726 8134
rect 11750 8132 11806 8134
rect 11510 7098 11566 7100
rect 11590 7098 11646 7100
rect 11670 7098 11726 7100
rect 11750 7098 11806 7100
rect 11510 7046 11556 7098
rect 11556 7046 11566 7098
rect 11590 7046 11620 7098
rect 11620 7046 11632 7098
rect 11632 7046 11646 7098
rect 11670 7046 11684 7098
rect 11684 7046 11696 7098
rect 11696 7046 11726 7098
rect 11750 7046 11760 7098
rect 11760 7046 11806 7098
rect 11510 7044 11566 7046
rect 11590 7044 11646 7046
rect 11670 7044 11726 7046
rect 11750 7044 11806 7046
rect 9659 5466 9715 5468
rect 9739 5466 9795 5468
rect 9819 5466 9875 5468
rect 9899 5466 9955 5468
rect 9659 5414 9705 5466
rect 9705 5414 9715 5466
rect 9739 5414 9769 5466
rect 9769 5414 9781 5466
rect 9781 5414 9795 5466
rect 9819 5414 9833 5466
rect 9833 5414 9845 5466
rect 9845 5414 9875 5466
rect 9899 5414 9909 5466
rect 9909 5414 9955 5466
rect 9659 5412 9715 5414
rect 9739 5412 9795 5414
rect 9819 5412 9875 5414
rect 9899 5412 9955 5414
rect 11510 6010 11566 6012
rect 11590 6010 11646 6012
rect 11670 6010 11726 6012
rect 11750 6010 11806 6012
rect 11510 5958 11556 6010
rect 11556 5958 11566 6010
rect 11590 5958 11620 6010
rect 11620 5958 11632 6010
rect 11632 5958 11646 6010
rect 11670 5958 11684 6010
rect 11684 5958 11696 6010
rect 11696 5958 11726 6010
rect 11750 5958 11760 6010
rect 11760 5958 11806 6010
rect 11510 5956 11566 5958
rect 11590 5956 11646 5958
rect 11670 5956 11726 5958
rect 11750 5956 11806 5958
rect 13361 15258 13417 15260
rect 13441 15258 13497 15260
rect 13521 15258 13577 15260
rect 13601 15258 13657 15260
rect 13361 15206 13407 15258
rect 13407 15206 13417 15258
rect 13441 15206 13471 15258
rect 13471 15206 13483 15258
rect 13483 15206 13497 15258
rect 13521 15206 13535 15258
rect 13535 15206 13547 15258
rect 13547 15206 13577 15258
rect 13601 15206 13611 15258
rect 13611 15206 13657 15258
rect 13361 15204 13417 15206
rect 13441 15204 13497 15206
rect 13521 15204 13577 15206
rect 13601 15204 13657 15206
rect 15212 14714 15268 14716
rect 15292 14714 15348 14716
rect 15372 14714 15428 14716
rect 15452 14714 15508 14716
rect 15212 14662 15258 14714
rect 15258 14662 15268 14714
rect 15292 14662 15322 14714
rect 15322 14662 15334 14714
rect 15334 14662 15348 14714
rect 15372 14662 15386 14714
rect 15386 14662 15398 14714
rect 15398 14662 15428 14714
rect 15452 14662 15462 14714
rect 15462 14662 15508 14714
rect 15212 14660 15268 14662
rect 15292 14660 15348 14662
rect 15372 14660 15428 14662
rect 15452 14660 15508 14662
rect 13361 14170 13417 14172
rect 13441 14170 13497 14172
rect 13521 14170 13577 14172
rect 13601 14170 13657 14172
rect 13361 14118 13407 14170
rect 13407 14118 13417 14170
rect 13441 14118 13471 14170
rect 13471 14118 13483 14170
rect 13483 14118 13497 14170
rect 13521 14118 13535 14170
rect 13535 14118 13547 14170
rect 13547 14118 13577 14170
rect 13601 14118 13611 14170
rect 13611 14118 13657 14170
rect 13361 14116 13417 14118
rect 13441 14116 13497 14118
rect 13521 14116 13577 14118
rect 13601 14116 13657 14118
rect 15014 13912 15070 13968
rect 15212 13626 15268 13628
rect 15292 13626 15348 13628
rect 15372 13626 15428 13628
rect 15452 13626 15508 13628
rect 15212 13574 15258 13626
rect 15258 13574 15268 13626
rect 15292 13574 15322 13626
rect 15322 13574 15334 13626
rect 15334 13574 15348 13626
rect 15372 13574 15386 13626
rect 15386 13574 15398 13626
rect 15398 13574 15428 13626
rect 15452 13574 15462 13626
rect 15462 13574 15508 13626
rect 15212 13572 15268 13574
rect 15292 13572 15348 13574
rect 15372 13572 15428 13574
rect 15452 13572 15508 13574
rect 15014 13132 15016 13152
rect 15016 13132 15068 13152
rect 15068 13132 15070 13152
rect 15014 13096 15070 13132
rect 13361 13082 13417 13084
rect 13441 13082 13497 13084
rect 13521 13082 13577 13084
rect 13601 13082 13657 13084
rect 13361 13030 13407 13082
rect 13407 13030 13417 13082
rect 13441 13030 13471 13082
rect 13471 13030 13483 13082
rect 13483 13030 13497 13082
rect 13521 13030 13535 13082
rect 13535 13030 13547 13082
rect 13547 13030 13577 13082
rect 13601 13030 13611 13082
rect 13611 13030 13657 13082
rect 13361 13028 13417 13030
rect 13441 13028 13497 13030
rect 13521 13028 13577 13030
rect 13601 13028 13657 13030
rect 15212 12538 15268 12540
rect 15292 12538 15348 12540
rect 15372 12538 15428 12540
rect 15452 12538 15508 12540
rect 15212 12486 15258 12538
rect 15258 12486 15268 12538
rect 15292 12486 15322 12538
rect 15322 12486 15334 12538
rect 15334 12486 15348 12538
rect 15372 12486 15386 12538
rect 15386 12486 15398 12538
rect 15398 12486 15428 12538
rect 15452 12486 15462 12538
rect 15462 12486 15508 12538
rect 15212 12484 15268 12486
rect 15292 12484 15348 12486
rect 15372 12484 15428 12486
rect 15452 12484 15508 12486
rect 15014 12280 15070 12336
rect 13361 11994 13417 11996
rect 13441 11994 13497 11996
rect 13521 11994 13577 11996
rect 13601 11994 13657 11996
rect 13361 11942 13407 11994
rect 13407 11942 13417 11994
rect 13441 11942 13471 11994
rect 13471 11942 13483 11994
rect 13483 11942 13497 11994
rect 13521 11942 13535 11994
rect 13535 11942 13547 11994
rect 13547 11942 13577 11994
rect 13601 11942 13611 11994
rect 13611 11942 13657 11994
rect 13361 11940 13417 11942
rect 13441 11940 13497 11942
rect 13521 11940 13577 11942
rect 13601 11940 13657 11942
rect 13361 10906 13417 10908
rect 13441 10906 13497 10908
rect 13521 10906 13577 10908
rect 13601 10906 13657 10908
rect 13361 10854 13407 10906
rect 13407 10854 13417 10906
rect 13441 10854 13471 10906
rect 13471 10854 13483 10906
rect 13483 10854 13497 10906
rect 13521 10854 13535 10906
rect 13535 10854 13547 10906
rect 13547 10854 13577 10906
rect 13601 10854 13611 10906
rect 13611 10854 13657 10906
rect 13361 10852 13417 10854
rect 13441 10852 13497 10854
rect 13521 10852 13577 10854
rect 13601 10852 13657 10854
rect 13361 9818 13417 9820
rect 13441 9818 13497 9820
rect 13521 9818 13577 9820
rect 13601 9818 13657 9820
rect 13361 9766 13407 9818
rect 13407 9766 13417 9818
rect 13441 9766 13471 9818
rect 13471 9766 13483 9818
rect 13483 9766 13497 9818
rect 13521 9766 13535 9818
rect 13535 9766 13547 9818
rect 13547 9766 13577 9818
rect 13601 9766 13611 9818
rect 13611 9766 13657 9818
rect 13361 9764 13417 9766
rect 13441 9764 13497 9766
rect 13521 9764 13577 9766
rect 13601 9764 13657 9766
rect 13361 8730 13417 8732
rect 13441 8730 13497 8732
rect 13521 8730 13577 8732
rect 13601 8730 13657 8732
rect 13361 8678 13407 8730
rect 13407 8678 13417 8730
rect 13441 8678 13471 8730
rect 13471 8678 13483 8730
rect 13483 8678 13497 8730
rect 13521 8678 13535 8730
rect 13535 8678 13547 8730
rect 13547 8678 13577 8730
rect 13601 8678 13611 8730
rect 13611 8678 13657 8730
rect 13361 8676 13417 8678
rect 13441 8676 13497 8678
rect 13521 8676 13577 8678
rect 13601 8676 13657 8678
rect 13726 7964 13728 7984
rect 13728 7964 13780 7984
rect 13780 7964 13782 7984
rect 13726 7928 13782 7964
rect 13361 7642 13417 7644
rect 13441 7642 13497 7644
rect 13521 7642 13577 7644
rect 13601 7642 13657 7644
rect 13361 7590 13407 7642
rect 13407 7590 13417 7642
rect 13441 7590 13471 7642
rect 13471 7590 13483 7642
rect 13483 7590 13497 7642
rect 13521 7590 13535 7642
rect 13535 7590 13547 7642
rect 13547 7590 13577 7642
rect 13601 7590 13611 7642
rect 13611 7590 13657 7642
rect 13361 7588 13417 7590
rect 13441 7588 13497 7590
rect 13521 7588 13577 7590
rect 13601 7588 13657 7590
rect 15658 11464 15714 11520
rect 15212 11450 15268 11452
rect 15292 11450 15348 11452
rect 15372 11450 15428 11452
rect 15452 11450 15508 11452
rect 15212 11398 15258 11450
rect 15258 11398 15268 11450
rect 15292 11398 15322 11450
rect 15322 11398 15334 11450
rect 15334 11398 15348 11450
rect 15372 11398 15386 11450
rect 15386 11398 15398 11450
rect 15398 11398 15428 11450
rect 15452 11398 15462 11450
rect 15462 11398 15508 11450
rect 15212 11396 15268 11398
rect 15292 11396 15348 11398
rect 15372 11396 15428 11398
rect 15452 11396 15508 11398
rect 14738 7384 14794 7440
rect 11886 5752 11942 5808
rect 13361 6554 13417 6556
rect 13441 6554 13497 6556
rect 13521 6554 13577 6556
rect 13601 6554 13657 6556
rect 13361 6502 13407 6554
rect 13407 6502 13417 6554
rect 13441 6502 13471 6554
rect 13471 6502 13483 6554
rect 13483 6502 13497 6554
rect 13521 6502 13535 6554
rect 13535 6502 13547 6554
rect 13547 6502 13577 6554
rect 13601 6502 13611 6554
rect 13611 6502 13657 6554
rect 13361 6500 13417 6502
rect 13441 6500 13497 6502
rect 13521 6500 13577 6502
rect 13601 6500 13657 6502
rect 13361 5466 13417 5468
rect 13441 5466 13497 5468
rect 13521 5466 13577 5468
rect 13601 5466 13657 5468
rect 13361 5414 13407 5466
rect 13407 5414 13417 5466
rect 13441 5414 13471 5466
rect 13471 5414 13483 5466
rect 13483 5414 13497 5466
rect 13521 5414 13535 5466
rect 13535 5414 13547 5466
rect 13547 5414 13577 5466
rect 13601 5414 13611 5466
rect 13611 5414 13657 5466
rect 13361 5412 13417 5414
rect 13441 5412 13497 5414
rect 13521 5412 13577 5414
rect 13601 5412 13657 5414
rect 15014 10668 15070 10704
rect 15014 10648 15016 10668
rect 15016 10648 15068 10668
rect 15068 10648 15070 10668
rect 15212 10362 15268 10364
rect 15292 10362 15348 10364
rect 15372 10362 15428 10364
rect 15452 10362 15508 10364
rect 15212 10310 15258 10362
rect 15258 10310 15268 10362
rect 15292 10310 15322 10362
rect 15322 10310 15334 10362
rect 15334 10310 15348 10362
rect 15372 10310 15386 10362
rect 15386 10310 15398 10362
rect 15398 10310 15428 10362
rect 15452 10310 15462 10362
rect 15462 10310 15508 10362
rect 15212 10308 15268 10310
rect 15292 10308 15348 10310
rect 15372 10308 15428 10310
rect 15452 10308 15508 10310
rect 15014 9868 15016 9888
rect 15016 9868 15068 9888
rect 15068 9868 15070 9888
rect 15014 9832 15070 9868
rect 15212 9274 15268 9276
rect 15292 9274 15348 9276
rect 15372 9274 15428 9276
rect 15452 9274 15508 9276
rect 15212 9222 15258 9274
rect 15258 9222 15268 9274
rect 15292 9222 15322 9274
rect 15322 9222 15334 9274
rect 15334 9222 15348 9274
rect 15372 9222 15386 9274
rect 15386 9222 15398 9274
rect 15398 9222 15428 9274
rect 15452 9222 15462 9274
rect 15462 9222 15508 9274
rect 15212 9220 15268 9222
rect 15292 9220 15348 9222
rect 15372 9220 15428 9222
rect 15452 9220 15508 9222
rect 15014 9016 15070 9072
rect 15212 8186 15268 8188
rect 15292 8186 15348 8188
rect 15372 8186 15428 8188
rect 15452 8186 15508 8188
rect 15212 8134 15258 8186
rect 15258 8134 15268 8186
rect 15292 8134 15322 8186
rect 15322 8134 15334 8186
rect 15334 8134 15348 8186
rect 15372 8134 15386 8186
rect 15386 8134 15398 8186
rect 15398 8134 15428 8186
rect 15452 8134 15462 8186
rect 15462 8134 15508 8186
rect 15212 8132 15268 8134
rect 15292 8132 15348 8134
rect 15372 8132 15428 8134
rect 15452 8132 15508 8134
rect 15212 7098 15268 7100
rect 15292 7098 15348 7100
rect 15372 7098 15428 7100
rect 15452 7098 15508 7100
rect 15212 7046 15258 7098
rect 15258 7046 15268 7098
rect 15292 7046 15322 7098
rect 15322 7046 15334 7098
rect 15334 7046 15348 7098
rect 15372 7046 15386 7098
rect 15386 7046 15398 7098
rect 15398 7046 15428 7098
rect 15452 7046 15462 7098
rect 15462 7046 15508 7098
rect 15212 7044 15268 7046
rect 15292 7044 15348 7046
rect 15372 7044 15428 7046
rect 15452 7044 15508 7046
rect 15014 6840 15070 6896
rect 14922 6568 14978 6624
rect 11510 4922 11566 4924
rect 11590 4922 11646 4924
rect 11670 4922 11726 4924
rect 11750 4922 11806 4924
rect 11510 4870 11556 4922
rect 11556 4870 11566 4922
rect 11590 4870 11620 4922
rect 11620 4870 11632 4922
rect 11632 4870 11646 4922
rect 11670 4870 11684 4922
rect 11684 4870 11696 4922
rect 11696 4870 11726 4922
rect 11750 4870 11760 4922
rect 11760 4870 11806 4922
rect 11510 4868 11566 4870
rect 11590 4868 11646 4870
rect 11670 4868 11726 4870
rect 11750 4868 11806 4870
rect 9659 4378 9715 4380
rect 9739 4378 9795 4380
rect 9819 4378 9875 4380
rect 9899 4378 9955 4380
rect 9659 4326 9705 4378
rect 9705 4326 9715 4378
rect 9739 4326 9769 4378
rect 9769 4326 9781 4378
rect 9781 4326 9795 4378
rect 9819 4326 9833 4378
rect 9833 4326 9845 4378
rect 9845 4326 9875 4378
rect 9899 4326 9909 4378
rect 9909 4326 9955 4378
rect 9659 4324 9715 4326
rect 9739 4324 9795 4326
rect 9819 4324 9875 4326
rect 9899 4324 9955 4326
rect 4106 2746 4162 2748
rect 4186 2746 4242 2748
rect 4266 2746 4322 2748
rect 4346 2746 4402 2748
rect 4106 2694 4152 2746
rect 4152 2694 4162 2746
rect 4186 2694 4216 2746
rect 4216 2694 4228 2746
rect 4228 2694 4242 2746
rect 4266 2694 4280 2746
rect 4280 2694 4292 2746
rect 4292 2694 4322 2746
rect 4346 2694 4356 2746
rect 4356 2694 4402 2746
rect 4106 2692 4162 2694
rect 4186 2692 4242 2694
rect 4266 2692 4322 2694
rect 4346 2692 4402 2694
rect 7808 2746 7864 2748
rect 7888 2746 7944 2748
rect 7968 2746 8024 2748
rect 8048 2746 8104 2748
rect 7808 2694 7854 2746
rect 7854 2694 7864 2746
rect 7888 2694 7918 2746
rect 7918 2694 7930 2746
rect 7930 2694 7944 2746
rect 7968 2694 7982 2746
rect 7982 2694 7994 2746
rect 7994 2694 8024 2746
rect 8048 2694 8058 2746
rect 8058 2694 8104 2746
rect 7808 2692 7864 2694
rect 7888 2692 7944 2694
rect 7968 2692 8024 2694
rect 8048 2692 8104 2694
rect 8298 2508 8354 2544
rect 8298 2488 8300 2508
rect 8300 2488 8352 2508
rect 8352 2488 8354 2508
rect 2255 2202 2311 2204
rect 2335 2202 2391 2204
rect 2415 2202 2471 2204
rect 2495 2202 2551 2204
rect 2255 2150 2301 2202
rect 2301 2150 2311 2202
rect 2335 2150 2365 2202
rect 2365 2150 2377 2202
rect 2377 2150 2391 2202
rect 2415 2150 2429 2202
rect 2429 2150 2441 2202
rect 2441 2150 2471 2202
rect 2495 2150 2505 2202
rect 2505 2150 2551 2202
rect 2255 2148 2311 2150
rect 2335 2148 2391 2150
rect 2415 2148 2471 2150
rect 2495 2148 2551 2150
rect 5957 2202 6013 2204
rect 6037 2202 6093 2204
rect 6117 2202 6173 2204
rect 6197 2202 6253 2204
rect 5957 2150 6003 2202
rect 6003 2150 6013 2202
rect 6037 2150 6067 2202
rect 6067 2150 6079 2202
rect 6079 2150 6093 2202
rect 6117 2150 6131 2202
rect 6131 2150 6143 2202
rect 6143 2150 6173 2202
rect 6197 2150 6207 2202
rect 6207 2150 6253 2202
rect 5957 2148 6013 2150
rect 6037 2148 6093 2150
rect 6117 2148 6173 2150
rect 6197 2148 6253 2150
rect 4106 1658 4162 1660
rect 4186 1658 4242 1660
rect 4266 1658 4322 1660
rect 4346 1658 4402 1660
rect 4106 1606 4152 1658
rect 4152 1606 4162 1658
rect 4186 1606 4216 1658
rect 4216 1606 4228 1658
rect 4228 1606 4242 1658
rect 4266 1606 4280 1658
rect 4280 1606 4292 1658
rect 4292 1606 4322 1658
rect 4346 1606 4356 1658
rect 4356 1606 4402 1658
rect 4106 1604 4162 1606
rect 4186 1604 4242 1606
rect 4266 1604 4322 1606
rect 4346 1604 4402 1606
rect 2255 1114 2311 1116
rect 2335 1114 2391 1116
rect 2415 1114 2471 1116
rect 2495 1114 2551 1116
rect 2255 1062 2301 1114
rect 2301 1062 2311 1114
rect 2335 1062 2365 1114
rect 2365 1062 2377 1114
rect 2377 1062 2391 1114
rect 2415 1062 2429 1114
rect 2429 1062 2441 1114
rect 2441 1062 2471 1114
rect 2495 1062 2505 1114
rect 2505 1062 2551 1114
rect 2255 1060 2311 1062
rect 2335 1060 2391 1062
rect 2415 1060 2471 1062
rect 2495 1060 2551 1062
rect 5957 1114 6013 1116
rect 6037 1114 6093 1116
rect 6117 1114 6173 1116
rect 6197 1114 6253 1116
rect 5957 1062 6003 1114
rect 6003 1062 6013 1114
rect 6037 1062 6067 1114
rect 6067 1062 6079 1114
rect 6079 1062 6093 1114
rect 6117 1062 6131 1114
rect 6131 1062 6143 1114
rect 6143 1062 6173 1114
rect 6197 1062 6207 1114
rect 6207 1062 6253 1114
rect 5957 1060 6013 1062
rect 6037 1060 6093 1062
rect 6117 1060 6173 1062
rect 6197 1060 6253 1062
rect 7808 1658 7864 1660
rect 7888 1658 7944 1660
rect 7968 1658 8024 1660
rect 8048 1658 8104 1660
rect 7808 1606 7854 1658
rect 7854 1606 7864 1658
rect 7888 1606 7918 1658
rect 7918 1606 7930 1658
rect 7930 1606 7944 1658
rect 7968 1606 7982 1658
rect 7982 1606 7994 1658
rect 7994 1606 8024 1658
rect 8048 1606 8058 1658
rect 8058 1606 8104 1658
rect 7808 1604 7864 1606
rect 7888 1604 7944 1606
rect 7968 1604 8024 1606
rect 8048 1604 8104 1606
rect 9659 3290 9715 3292
rect 9739 3290 9795 3292
rect 9819 3290 9875 3292
rect 9899 3290 9955 3292
rect 9659 3238 9705 3290
rect 9705 3238 9715 3290
rect 9739 3238 9769 3290
rect 9769 3238 9781 3290
rect 9781 3238 9795 3290
rect 9819 3238 9833 3290
rect 9833 3238 9845 3290
rect 9845 3238 9875 3290
rect 9899 3238 9909 3290
rect 9909 3238 9955 3290
rect 9659 3236 9715 3238
rect 9739 3236 9795 3238
rect 9819 3236 9875 3238
rect 9899 3236 9955 3238
rect 9659 2202 9715 2204
rect 9739 2202 9795 2204
rect 9819 2202 9875 2204
rect 9899 2202 9955 2204
rect 9659 2150 9705 2202
rect 9705 2150 9715 2202
rect 9739 2150 9769 2202
rect 9769 2150 9781 2202
rect 9781 2150 9795 2202
rect 9819 2150 9833 2202
rect 9833 2150 9845 2202
rect 9845 2150 9875 2202
rect 9899 2150 9909 2202
rect 9909 2150 9955 2202
rect 9659 2148 9715 2150
rect 9739 2148 9795 2150
rect 9819 2148 9875 2150
rect 9899 2148 9955 2150
rect 10046 1828 10102 1864
rect 10046 1808 10048 1828
rect 10048 1808 10100 1828
rect 10100 1808 10102 1828
rect 9659 1114 9715 1116
rect 9739 1114 9795 1116
rect 9819 1114 9875 1116
rect 9899 1114 9955 1116
rect 9659 1062 9705 1114
rect 9705 1062 9715 1114
rect 9739 1062 9769 1114
rect 9769 1062 9781 1114
rect 9781 1062 9795 1114
rect 9819 1062 9833 1114
rect 9833 1062 9845 1114
rect 9845 1062 9875 1114
rect 9899 1062 9909 1114
rect 9909 1062 9955 1114
rect 9659 1060 9715 1062
rect 9739 1060 9795 1062
rect 9819 1060 9875 1062
rect 9899 1060 9955 1062
rect 11510 3834 11566 3836
rect 11590 3834 11646 3836
rect 11670 3834 11726 3836
rect 11750 3834 11806 3836
rect 11510 3782 11556 3834
rect 11556 3782 11566 3834
rect 11590 3782 11620 3834
rect 11620 3782 11632 3834
rect 11632 3782 11646 3834
rect 11670 3782 11684 3834
rect 11684 3782 11696 3834
rect 11696 3782 11726 3834
rect 11750 3782 11760 3834
rect 11760 3782 11806 3834
rect 11510 3780 11566 3782
rect 11590 3780 11646 3782
rect 11670 3780 11726 3782
rect 11750 3780 11806 3782
rect 13082 4120 13138 4176
rect 13361 4378 13417 4380
rect 13441 4378 13497 4380
rect 13521 4378 13577 4380
rect 13601 4378 13657 4380
rect 13361 4326 13407 4378
rect 13407 4326 13417 4378
rect 13441 4326 13471 4378
rect 13471 4326 13483 4378
rect 13483 4326 13497 4378
rect 13521 4326 13535 4378
rect 13535 4326 13547 4378
rect 13547 4326 13577 4378
rect 13601 4326 13611 4378
rect 13611 4326 13657 4378
rect 13361 4324 13417 4326
rect 13441 4324 13497 4326
rect 13521 4324 13577 4326
rect 13601 4324 13657 4326
rect 15212 6010 15268 6012
rect 15292 6010 15348 6012
rect 15372 6010 15428 6012
rect 15452 6010 15508 6012
rect 15212 5958 15258 6010
rect 15258 5958 15268 6010
rect 15292 5958 15322 6010
rect 15322 5958 15334 6010
rect 15334 5958 15348 6010
rect 15372 5958 15386 6010
rect 15386 5958 15398 6010
rect 15398 5958 15428 6010
rect 15452 5958 15462 6010
rect 15462 5958 15508 6010
rect 15212 5956 15268 5958
rect 15292 5956 15348 5958
rect 15372 5956 15428 5958
rect 15452 5956 15508 5958
rect 13910 5788 13912 5808
rect 13912 5788 13964 5808
rect 13964 5788 13966 5808
rect 13910 5752 13966 5788
rect 13910 4120 13966 4176
rect 11510 2746 11566 2748
rect 11590 2746 11646 2748
rect 11670 2746 11726 2748
rect 11750 2746 11806 2748
rect 11510 2694 11556 2746
rect 11556 2694 11566 2746
rect 11590 2694 11620 2746
rect 11620 2694 11632 2746
rect 11632 2694 11646 2746
rect 11670 2694 11684 2746
rect 11684 2694 11696 2746
rect 11696 2694 11726 2746
rect 11750 2694 11760 2746
rect 11760 2694 11806 2746
rect 11510 2692 11566 2694
rect 11590 2692 11646 2694
rect 11670 2692 11726 2694
rect 11750 2692 11806 2694
rect 11510 1658 11566 1660
rect 11590 1658 11646 1660
rect 11670 1658 11726 1660
rect 11750 1658 11806 1660
rect 11510 1606 11556 1658
rect 11556 1606 11566 1658
rect 11590 1606 11620 1658
rect 11620 1606 11632 1658
rect 11632 1606 11646 1658
rect 11670 1606 11684 1658
rect 11684 1606 11696 1658
rect 11696 1606 11726 1658
rect 11750 1606 11760 1658
rect 11760 1606 11806 1658
rect 11510 1604 11566 1606
rect 11590 1604 11646 1606
rect 11670 1604 11726 1606
rect 11750 1604 11806 1606
rect 13361 3290 13417 3292
rect 13441 3290 13497 3292
rect 13521 3290 13577 3292
rect 13601 3290 13657 3292
rect 13361 3238 13407 3290
rect 13407 3238 13417 3290
rect 13441 3238 13471 3290
rect 13471 3238 13483 3290
rect 13483 3238 13497 3290
rect 13521 3238 13535 3290
rect 13535 3238 13547 3290
rect 13547 3238 13577 3290
rect 13601 3238 13611 3290
rect 13611 3238 13657 3290
rect 13361 3236 13417 3238
rect 13441 3236 13497 3238
rect 13521 3236 13577 3238
rect 13601 3236 13657 3238
rect 13361 2202 13417 2204
rect 13441 2202 13497 2204
rect 13521 2202 13577 2204
rect 13601 2202 13657 2204
rect 13361 2150 13407 2202
rect 13407 2150 13417 2202
rect 13441 2150 13471 2202
rect 13471 2150 13483 2202
rect 13483 2150 13497 2202
rect 13521 2150 13535 2202
rect 13535 2150 13547 2202
rect 13547 2150 13577 2202
rect 13601 2150 13611 2202
rect 13611 2150 13657 2202
rect 13361 2148 13417 2150
rect 13441 2148 13497 2150
rect 13521 2148 13577 2150
rect 13601 2148 13657 2150
rect 15658 8200 15714 8256
rect 15934 6840 15990 6896
rect 15566 5752 15622 5808
rect 15934 4936 15990 4992
rect 15212 4922 15268 4924
rect 15292 4922 15348 4924
rect 15372 4922 15428 4924
rect 15452 4922 15508 4924
rect 15212 4870 15258 4922
rect 15258 4870 15268 4922
rect 15292 4870 15322 4922
rect 15322 4870 15334 4922
rect 15334 4870 15348 4922
rect 15372 4870 15386 4922
rect 15386 4870 15398 4922
rect 15398 4870 15428 4922
rect 15452 4870 15462 4922
rect 15462 4870 15508 4922
rect 15212 4868 15268 4870
rect 15292 4868 15348 4870
rect 15372 4868 15428 4870
rect 15452 4868 15508 4870
rect 15014 4120 15070 4176
rect 15212 3834 15268 3836
rect 15292 3834 15348 3836
rect 15372 3834 15428 3836
rect 15452 3834 15508 3836
rect 15212 3782 15258 3834
rect 15258 3782 15268 3834
rect 15292 3782 15322 3834
rect 15322 3782 15334 3834
rect 15334 3782 15348 3834
rect 15372 3782 15386 3834
rect 15386 3782 15398 3834
rect 15398 3782 15428 3834
rect 15452 3782 15462 3834
rect 15462 3782 15508 3834
rect 15212 3780 15268 3782
rect 15292 3780 15348 3782
rect 15372 3780 15428 3782
rect 15452 3780 15508 3782
rect 15014 3304 15070 3360
rect 15212 2746 15268 2748
rect 15292 2746 15348 2748
rect 15372 2746 15428 2748
rect 15452 2746 15508 2748
rect 15212 2694 15258 2746
rect 15258 2694 15268 2746
rect 15292 2694 15322 2746
rect 15322 2694 15334 2746
rect 15334 2694 15348 2746
rect 15372 2694 15386 2746
rect 15386 2694 15398 2746
rect 15398 2694 15428 2746
rect 15452 2694 15462 2746
rect 15462 2694 15508 2746
rect 15212 2692 15268 2694
rect 15292 2692 15348 2694
rect 15372 2692 15428 2694
rect 15452 2692 15508 2694
rect 15014 2508 15070 2544
rect 15014 2488 15016 2508
rect 15016 2488 15068 2508
rect 15068 2488 15070 2508
rect 15014 1808 15070 1864
rect 15658 1672 15714 1728
rect 15212 1658 15268 1660
rect 15292 1658 15348 1660
rect 15372 1658 15428 1660
rect 15452 1658 15508 1660
rect 15212 1606 15258 1658
rect 15258 1606 15268 1658
rect 15292 1606 15322 1658
rect 15322 1606 15334 1658
rect 15334 1606 15348 1658
rect 15372 1606 15386 1658
rect 15386 1606 15398 1658
rect 15398 1606 15428 1658
rect 15452 1606 15462 1658
rect 15462 1606 15508 1658
rect 15212 1604 15268 1606
rect 15292 1604 15348 1606
rect 15372 1604 15428 1606
rect 15452 1604 15508 1606
rect 13361 1114 13417 1116
rect 13441 1114 13497 1116
rect 13521 1114 13577 1116
rect 13601 1114 13657 1116
rect 13361 1062 13407 1114
rect 13407 1062 13417 1114
rect 13441 1062 13471 1114
rect 13471 1062 13483 1114
rect 13483 1062 13497 1114
rect 13521 1062 13535 1114
rect 13535 1062 13547 1114
rect 13547 1062 13577 1114
rect 13601 1062 13611 1114
rect 13611 1062 13657 1114
rect 13361 1060 13417 1062
rect 13441 1060 13497 1062
rect 13521 1060 13577 1062
rect 13601 1060 13657 1062
rect 4106 570 4162 572
rect 4186 570 4242 572
rect 4266 570 4322 572
rect 4346 570 4402 572
rect 4106 518 4152 570
rect 4152 518 4162 570
rect 4186 518 4216 570
rect 4216 518 4228 570
rect 4228 518 4242 570
rect 4266 518 4280 570
rect 4280 518 4292 570
rect 4292 518 4322 570
rect 4346 518 4356 570
rect 4356 518 4402 570
rect 4106 516 4162 518
rect 4186 516 4242 518
rect 4266 516 4322 518
rect 4346 516 4402 518
rect 7808 570 7864 572
rect 7888 570 7944 572
rect 7968 570 8024 572
rect 8048 570 8104 572
rect 7808 518 7854 570
rect 7854 518 7864 570
rect 7888 518 7918 570
rect 7918 518 7930 570
rect 7930 518 7944 570
rect 7968 518 7982 570
rect 7982 518 7994 570
rect 7994 518 8024 570
rect 8048 518 8058 570
rect 8058 518 8104 570
rect 7808 516 7864 518
rect 7888 516 7944 518
rect 7968 516 8024 518
rect 8048 516 8104 518
rect 11510 570 11566 572
rect 11590 570 11646 572
rect 11670 570 11726 572
rect 11750 570 11806 572
rect 11510 518 11556 570
rect 11556 518 11566 570
rect 11590 518 11620 570
rect 11620 518 11632 570
rect 11632 518 11646 570
rect 11670 518 11684 570
rect 11684 518 11696 570
rect 11696 518 11726 570
rect 11750 518 11760 570
rect 11760 518 11806 570
rect 11510 516 11566 518
rect 11590 516 11646 518
rect 11670 516 11726 518
rect 11750 516 11806 518
rect 15212 570 15268 572
rect 15292 570 15348 572
rect 15372 570 15428 572
rect 15452 570 15508 572
rect 15212 518 15258 570
rect 15258 518 15268 570
rect 15292 518 15322 570
rect 15322 518 15334 570
rect 15334 518 15348 570
rect 15372 518 15386 570
rect 15386 518 15398 570
rect 15398 518 15428 570
rect 15452 518 15462 570
rect 15462 518 15508 570
rect 15212 516 15268 518
rect 15292 516 15348 518
rect 15372 516 15428 518
rect 15452 516 15508 518
<< metal3 >>
rect 2245 15264 2561 15265
rect 2245 15200 2251 15264
rect 2315 15200 2331 15264
rect 2395 15200 2411 15264
rect 2475 15200 2491 15264
rect 2555 15200 2561 15264
rect 2245 15199 2561 15200
rect 5947 15264 6263 15265
rect 5947 15200 5953 15264
rect 6017 15200 6033 15264
rect 6097 15200 6113 15264
rect 6177 15200 6193 15264
rect 6257 15200 6263 15264
rect 5947 15199 6263 15200
rect 9649 15264 9965 15265
rect 9649 15200 9655 15264
rect 9719 15200 9735 15264
rect 9799 15200 9815 15264
rect 9879 15200 9895 15264
rect 9959 15200 9965 15264
rect 9649 15199 9965 15200
rect 13351 15264 13667 15265
rect 13351 15200 13357 15264
rect 13421 15200 13437 15264
rect 13501 15200 13517 15264
rect 13581 15200 13597 15264
rect 13661 15200 13667 15264
rect 13351 15199 13667 15200
rect 4096 14720 4412 14721
rect 4096 14656 4102 14720
rect 4166 14656 4182 14720
rect 4246 14656 4262 14720
rect 4326 14656 4342 14720
rect 4406 14656 4412 14720
rect 4096 14655 4412 14656
rect 7798 14720 8114 14721
rect 7798 14656 7804 14720
rect 7868 14656 7884 14720
rect 7948 14656 7964 14720
rect 8028 14656 8044 14720
rect 8108 14656 8114 14720
rect 7798 14655 8114 14656
rect 11500 14720 11816 14721
rect 11500 14656 11506 14720
rect 11570 14656 11586 14720
rect 11650 14656 11666 14720
rect 11730 14656 11746 14720
rect 11810 14656 11816 14720
rect 11500 14655 11816 14656
rect 15202 14720 15518 14721
rect 15202 14656 15208 14720
rect 15272 14656 15288 14720
rect 15352 14656 15368 14720
rect 15432 14656 15448 14720
rect 15512 14656 15518 14720
rect 15202 14655 15518 14656
rect 2245 14176 2561 14177
rect 2245 14112 2251 14176
rect 2315 14112 2331 14176
rect 2395 14112 2411 14176
rect 2475 14112 2491 14176
rect 2555 14112 2561 14176
rect 2245 14111 2561 14112
rect 5947 14176 6263 14177
rect 5947 14112 5953 14176
rect 6017 14112 6033 14176
rect 6097 14112 6113 14176
rect 6177 14112 6193 14176
rect 6257 14112 6263 14176
rect 5947 14111 6263 14112
rect 9649 14176 9965 14177
rect 9649 14112 9655 14176
rect 9719 14112 9735 14176
rect 9799 14112 9815 14176
rect 9879 14112 9895 14176
rect 9959 14112 9965 14176
rect 9649 14111 9965 14112
rect 13351 14176 13667 14177
rect 13351 14112 13357 14176
rect 13421 14112 13437 14176
rect 13501 14112 13517 14176
rect 13581 14112 13597 14176
rect 13661 14112 13667 14176
rect 13351 14111 13667 14112
rect 15009 13970 15075 13973
rect 15600 13970 16000 14000
rect 15009 13968 16000 13970
rect 15009 13912 15014 13968
rect 15070 13912 16000 13968
rect 15009 13910 16000 13912
rect 15009 13907 15075 13910
rect 15600 13880 16000 13910
rect 4096 13632 4412 13633
rect 4096 13568 4102 13632
rect 4166 13568 4182 13632
rect 4246 13568 4262 13632
rect 4326 13568 4342 13632
rect 4406 13568 4412 13632
rect 4096 13567 4412 13568
rect 7798 13632 8114 13633
rect 7798 13568 7804 13632
rect 7868 13568 7884 13632
rect 7948 13568 7964 13632
rect 8028 13568 8044 13632
rect 8108 13568 8114 13632
rect 7798 13567 8114 13568
rect 11500 13632 11816 13633
rect 11500 13568 11506 13632
rect 11570 13568 11586 13632
rect 11650 13568 11666 13632
rect 11730 13568 11746 13632
rect 11810 13568 11816 13632
rect 11500 13567 11816 13568
rect 15202 13632 15518 13633
rect 15202 13568 15208 13632
rect 15272 13568 15288 13632
rect 15352 13568 15368 13632
rect 15432 13568 15448 13632
rect 15512 13568 15518 13632
rect 15202 13567 15518 13568
rect 15009 13154 15075 13157
rect 15600 13154 16000 13184
rect 15009 13152 16000 13154
rect 15009 13096 15014 13152
rect 15070 13096 16000 13152
rect 15009 13094 16000 13096
rect 15009 13091 15075 13094
rect 2245 13088 2561 13089
rect 2245 13024 2251 13088
rect 2315 13024 2331 13088
rect 2395 13024 2411 13088
rect 2475 13024 2491 13088
rect 2555 13024 2561 13088
rect 2245 13023 2561 13024
rect 5947 13088 6263 13089
rect 5947 13024 5953 13088
rect 6017 13024 6033 13088
rect 6097 13024 6113 13088
rect 6177 13024 6193 13088
rect 6257 13024 6263 13088
rect 5947 13023 6263 13024
rect 9649 13088 9965 13089
rect 9649 13024 9655 13088
rect 9719 13024 9735 13088
rect 9799 13024 9815 13088
rect 9879 13024 9895 13088
rect 9959 13024 9965 13088
rect 9649 13023 9965 13024
rect 13351 13088 13667 13089
rect 13351 13024 13357 13088
rect 13421 13024 13437 13088
rect 13501 13024 13517 13088
rect 13581 13024 13597 13088
rect 13661 13024 13667 13088
rect 15600 13064 16000 13094
rect 13351 13023 13667 13024
rect 4096 12544 4412 12545
rect 4096 12480 4102 12544
rect 4166 12480 4182 12544
rect 4246 12480 4262 12544
rect 4326 12480 4342 12544
rect 4406 12480 4412 12544
rect 4096 12479 4412 12480
rect 7798 12544 8114 12545
rect 7798 12480 7804 12544
rect 7868 12480 7884 12544
rect 7948 12480 7964 12544
rect 8028 12480 8044 12544
rect 8108 12480 8114 12544
rect 7798 12479 8114 12480
rect 11500 12544 11816 12545
rect 11500 12480 11506 12544
rect 11570 12480 11586 12544
rect 11650 12480 11666 12544
rect 11730 12480 11746 12544
rect 11810 12480 11816 12544
rect 11500 12479 11816 12480
rect 15202 12544 15518 12545
rect 15202 12480 15208 12544
rect 15272 12480 15288 12544
rect 15352 12480 15368 12544
rect 15432 12480 15448 12544
rect 15512 12480 15518 12544
rect 15202 12479 15518 12480
rect 15009 12338 15075 12341
rect 15600 12338 16000 12368
rect 15009 12336 16000 12338
rect 15009 12280 15014 12336
rect 15070 12280 16000 12336
rect 15009 12278 16000 12280
rect 15009 12275 15075 12278
rect 15600 12248 16000 12278
rect 2245 12000 2561 12001
rect 2245 11936 2251 12000
rect 2315 11936 2331 12000
rect 2395 11936 2411 12000
rect 2475 11936 2491 12000
rect 2555 11936 2561 12000
rect 2245 11935 2561 11936
rect 5947 12000 6263 12001
rect 5947 11936 5953 12000
rect 6017 11936 6033 12000
rect 6097 11936 6113 12000
rect 6177 11936 6193 12000
rect 6257 11936 6263 12000
rect 5947 11935 6263 11936
rect 9649 12000 9965 12001
rect 9649 11936 9655 12000
rect 9719 11936 9735 12000
rect 9799 11936 9815 12000
rect 9879 11936 9895 12000
rect 9959 11936 9965 12000
rect 9649 11935 9965 11936
rect 13351 12000 13667 12001
rect 13351 11936 13357 12000
rect 13421 11936 13437 12000
rect 13501 11936 13517 12000
rect 13581 11936 13597 12000
rect 13661 11936 13667 12000
rect 13351 11935 13667 11936
rect 15600 11520 16000 11552
rect 15600 11464 15658 11520
rect 15714 11464 16000 11520
rect 4096 11456 4412 11457
rect 4096 11392 4102 11456
rect 4166 11392 4182 11456
rect 4246 11392 4262 11456
rect 4326 11392 4342 11456
rect 4406 11392 4412 11456
rect 4096 11391 4412 11392
rect 7798 11456 8114 11457
rect 7798 11392 7804 11456
rect 7868 11392 7884 11456
rect 7948 11392 7964 11456
rect 8028 11392 8044 11456
rect 8108 11392 8114 11456
rect 7798 11391 8114 11392
rect 11500 11456 11816 11457
rect 11500 11392 11506 11456
rect 11570 11392 11586 11456
rect 11650 11392 11666 11456
rect 11730 11392 11746 11456
rect 11810 11392 11816 11456
rect 11500 11391 11816 11392
rect 15202 11456 15518 11457
rect 15202 11392 15208 11456
rect 15272 11392 15288 11456
rect 15352 11392 15368 11456
rect 15432 11392 15448 11456
rect 15512 11392 15518 11456
rect 15600 11432 16000 11464
rect 15202 11391 15518 11392
rect 2245 10912 2561 10913
rect 2245 10848 2251 10912
rect 2315 10848 2331 10912
rect 2395 10848 2411 10912
rect 2475 10848 2491 10912
rect 2555 10848 2561 10912
rect 2245 10847 2561 10848
rect 5947 10912 6263 10913
rect 5947 10848 5953 10912
rect 6017 10848 6033 10912
rect 6097 10848 6113 10912
rect 6177 10848 6193 10912
rect 6257 10848 6263 10912
rect 5947 10847 6263 10848
rect 9649 10912 9965 10913
rect 9649 10848 9655 10912
rect 9719 10848 9735 10912
rect 9799 10848 9815 10912
rect 9879 10848 9895 10912
rect 9959 10848 9965 10912
rect 9649 10847 9965 10848
rect 13351 10912 13667 10913
rect 13351 10848 13357 10912
rect 13421 10848 13437 10912
rect 13501 10848 13517 10912
rect 13581 10848 13597 10912
rect 13661 10848 13667 10912
rect 13351 10847 13667 10848
rect 15009 10706 15075 10709
rect 15600 10706 16000 10736
rect 15009 10704 16000 10706
rect 15009 10648 15014 10704
rect 15070 10648 16000 10704
rect 15009 10646 16000 10648
rect 15009 10643 15075 10646
rect 15600 10616 16000 10646
rect 4096 10368 4412 10369
rect 4096 10304 4102 10368
rect 4166 10304 4182 10368
rect 4246 10304 4262 10368
rect 4326 10304 4342 10368
rect 4406 10304 4412 10368
rect 4096 10303 4412 10304
rect 7798 10368 8114 10369
rect 7798 10304 7804 10368
rect 7868 10304 7884 10368
rect 7948 10304 7964 10368
rect 8028 10304 8044 10368
rect 8108 10304 8114 10368
rect 7798 10303 8114 10304
rect 11500 10368 11816 10369
rect 11500 10304 11506 10368
rect 11570 10304 11586 10368
rect 11650 10304 11666 10368
rect 11730 10304 11746 10368
rect 11810 10304 11816 10368
rect 11500 10303 11816 10304
rect 15202 10368 15518 10369
rect 15202 10304 15208 10368
rect 15272 10304 15288 10368
rect 15352 10304 15368 10368
rect 15432 10304 15448 10368
rect 15512 10304 15518 10368
rect 15202 10303 15518 10304
rect 15009 9890 15075 9893
rect 15600 9890 16000 9920
rect 15009 9888 16000 9890
rect 15009 9832 15014 9888
rect 15070 9832 16000 9888
rect 15009 9830 16000 9832
rect 15009 9827 15075 9830
rect 2245 9824 2561 9825
rect 2245 9760 2251 9824
rect 2315 9760 2331 9824
rect 2395 9760 2411 9824
rect 2475 9760 2491 9824
rect 2555 9760 2561 9824
rect 2245 9759 2561 9760
rect 5947 9824 6263 9825
rect 5947 9760 5953 9824
rect 6017 9760 6033 9824
rect 6097 9760 6113 9824
rect 6177 9760 6193 9824
rect 6257 9760 6263 9824
rect 5947 9759 6263 9760
rect 9649 9824 9965 9825
rect 9649 9760 9655 9824
rect 9719 9760 9735 9824
rect 9799 9760 9815 9824
rect 9879 9760 9895 9824
rect 9959 9760 9965 9824
rect 9649 9759 9965 9760
rect 13351 9824 13667 9825
rect 13351 9760 13357 9824
rect 13421 9760 13437 9824
rect 13501 9760 13517 9824
rect 13581 9760 13597 9824
rect 13661 9760 13667 9824
rect 15600 9800 16000 9830
rect 13351 9759 13667 9760
rect 4096 9280 4412 9281
rect 4096 9216 4102 9280
rect 4166 9216 4182 9280
rect 4246 9216 4262 9280
rect 4326 9216 4342 9280
rect 4406 9216 4412 9280
rect 4096 9215 4412 9216
rect 7798 9280 8114 9281
rect 7798 9216 7804 9280
rect 7868 9216 7884 9280
rect 7948 9216 7964 9280
rect 8028 9216 8044 9280
rect 8108 9216 8114 9280
rect 7798 9215 8114 9216
rect 11500 9280 11816 9281
rect 11500 9216 11506 9280
rect 11570 9216 11586 9280
rect 11650 9216 11666 9280
rect 11730 9216 11746 9280
rect 11810 9216 11816 9280
rect 11500 9215 11816 9216
rect 15202 9280 15518 9281
rect 15202 9216 15208 9280
rect 15272 9216 15288 9280
rect 15352 9216 15368 9280
rect 15432 9216 15448 9280
rect 15512 9216 15518 9280
rect 15202 9215 15518 9216
rect 9765 9074 9831 9077
rect 10501 9074 10567 9077
rect 9765 9072 10567 9074
rect 9765 9016 9770 9072
rect 9826 9016 10506 9072
rect 10562 9016 10567 9072
rect 9765 9014 10567 9016
rect 9765 9011 9831 9014
rect 10501 9011 10567 9014
rect 15009 9074 15075 9077
rect 15600 9074 16000 9104
rect 15009 9072 16000 9074
rect 15009 9016 15014 9072
rect 15070 9016 16000 9072
rect 15009 9014 16000 9016
rect 15009 9011 15075 9014
rect 15600 8984 16000 9014
rect 2245 8736 2561 8737
rect 2245 8672 2251 8736
rect 2315 8672 2331 8736
rect 2395 8672 2411 8736
rect 2475 8672 2491 8736
rect 2555 8672 2561 8736
rect 2245 8671 2561 8672
rect 5947 8736 6263 8737
rect 5947 8672 5953 8736
rect 6017 8672 6033 8736
rect 6097 8672 6113 8736
rect 6177 8672 6193 8736
rect 6257 8672 6263 8736
rect 5947 8671 6263 8672
rect 9649 8736 9965 8737
rect 9649 8672 9655 8736
rect 9719 8672 9735 8736
rect 9799 8672 9815 8736
rect 9879 8672 9895 8736
rect 9959 8672 9965 8736
rect 9649 8671 9965 8672
rect 13351 8736 13667 8737
rect 13351 8672 13357 8736
rect 13421 8672 13437 8736
rect 13501 8672 13517 8736
rect 13581 8672 13597 8736
rect 13661 8672 13667 8736
rect 13351 8671 13667 8672
rect 15600 8256 16000 8288
rect 15600 8200 15658 8256
rect 15714 8200 16000 8256
rect 4096 8192 4412 8193
rect 4096 8128 4102 8192
rect 4166 8128 4182 8192
rect 4246 8128 4262 8192
rect 4326 8128 4342 8192
rect 4406 8128 4412 8192
rect 4096 8127 4412 8128
rect 7798 8192 8114 8193
rect 7798 8128 7804 8192
rect 7868 8128 7884 8192
rect 7948 8128 7964 8192
rect 8028 8128 8044 8192
rect 8108 8128 8114 8192
rect 7798 8127 8114 8128
rect 11500 8192 11816 8193
rect 11500 8128 11506 8192
rect 11570 8128 11586 8192
rect 11650 8128 11666 8192
rect 11730 8128 11746 8192
rect 11810 8128 11816 8192
rect 11500 8127 11816 8128
rect 15202 8192 15518 8193
rect 15202 8128 15208 8192
rect 15272 8128 15288 8192
rect 15352 8128 15368 8192
rect 15432 8128 15448 8192
rect 15512 8128 15518 8192
rect 15600 8168 16000 8200
rect 15202 8127 15518 8128
rect 9213 7986 9279 7989
rect 13721 7986 13787 7989
rect 9213 7984 13787 7986
rect 9213 7928 9218 7984
rect 9274 7928 13726 7984
rect 13782 7928 13787 7984
rect 9213 7926 13787 7928
rect 9213 7923 9279 7926
rect 13721 7923 13787 7926
rect 2245 7648 2561 7649
rect 2245 7584 2251 7648
rect 2315 7584 2331 7648
rect 2395 7584 2411 7648
rect 2475 7584 2491 7648
rect 2555 7584 2561 7648
rect 2245 7583 2561 7584
rect 5947 7648 6263 7649
rect 5947 7584 5953 7648
rect 6017 7584 6033 7648
rect 6097 7584 6113 7648
rect 6177 7584 6193 7648
rect 6257 7584 6263 7648
rect 5947 7583 6263 7584
rect 9649 7648 9965 7649
rect 9649 7584 9655 7648
rect 9719 7584 9735 7648
rect 9799 7584 9815 7648
rect 9879 7584 9895 7648
rect 9959 7584 9965 7648
rect 9649 7583 9965 7584
rect 13351 7648 13667 7649
rect 13351 7584 13357 7648
rect 13421 7584 13437 7648
rect 13501 7584 13517 7648
rect 13581 7584 13597 7648
rect 13661 7584 13667 7648
rect 13351 7583 13667 7584
rect 14733 7442 14799 7445
rect 15600 7442 16000 7472
rect 14733 7440 16000 7442
rect 14733 7384 14738 7440
rect 14794 7384 16000 7440
rect 14733 7382 16000 7384
rect 14733 7379 14799 7382
rect 15600 7352 16000 7382
rect 4096 7104 4412 7105
rect 4096 7040 4102 7104
rect 4166 7040 4182 7104
rect 4246 7040 4262 7104
rect 4326 7040 4342 7104
rect 4406 7040 4412 7104
rect 4096 7039 4412 7040
rect 7798 7104 8114 7105
rect 7798 7040 7804 7104
rect 7868 7040 7884 7104
rect 7948 7040 7964 7104
rect 8028 7040 8044 7104
rect 8108 7040 8114 7104
rect 7798 7039 8114 7040
rect 11500 7104 11816 7105
rect 11500 7040 11506 7104
rect 11570 7040 11586 7104
rect 11650 7040 11666 7104
rect 11730 7040 11746 7104
rect 11810 7040 11816 7104
rect 11500 7039 11816 7040
rect 15202 7104 15518 7105
rect 15202 7040 15208 7104
rect 15272 7040 15288 7104
rect 15352 7040 15368 7104
rect 15432 7040 15448 7104
rect 15512 7040 15518 7104
rect 15202 7039 15518 7040
rect 9213 6898 9279 6901
rect 15009 6898 15075 6901
rect 15929 6898 15995 6901
rect 9213 6896 15995 6898
rect 9213 6840 9218 6896
rect 9274 6840 15014 6896
rect 15070 6840 15934 6896
rect 15990 6840 15995 6896
rect 9213 6838 15995 6840
rect 9213 6835 9279 6838
rect 15009 6835 15075 6838
rect 15929 6835 15995 6838
rect 14917 6626 14983 6629
rect 15600 6626 16000 6656
rect 14917 6624 16000 6626
rect 14917 6568 14922 6624
rect 14978 6568 16000 6624
rect 14917 6566 16000 6568
rect 14917 6563 14983 6566
rect 2245 6560 2561 6561
rect 2245 6496 2251 6560
rect 2315 6496 2331 6560
rect 2395 6496 2411 6560
rect 2475 6496 2491 6560
rect 2555 6496 2561 6560
rect 2245 6495 2561 6496
rect 5947 6560 6263 6561
rect 5947 6496 5953 6560
rect 6017 6496 6033 6560
rect 6097 6496 6113 6560
rect 6177 6496 6193 6560
rect 6257 6496 6263 6560
rect 5947 6495 6263 6496
rect 9649 6560 9965 6561
rect 9649 6496 9655 6560
rect 9719 6496 9735 6560
rect 9799 6496 9815 6560
rect 9879 6496 9895 6560
rect 9959 6496 9965 6560
rect 9649 6495 9965 6496
rect 13351 6560 13667 6561
rect 13351 6496 13357 6560
rect 13421 6496 13437 6560
rect 13501 6496 13517 6560
rect 13581 6496 13597 6560
rect 13661 6496 13667 6560
rect 15600 6536 16000 6566
rect 13351 6495 13667 6496
rect 4096 6016 4412 6017
rect 4096 5952 4102 6016
rect 4166 5952 4182 6016
rect 4246 5952 4262 6016
rect 4326 5952 4342 6016
rect 4406 5952 4412 6016
rect 4096 5951 4412 5952
rect 7798 6016 8114 6017
rect 7798 5952 7804 6016
rect 7868 5952 7884 6016
rect 7948 5952 7964 6016
rect 8028 5952 8044 6016
rect 8108 5952 8114 6016
rect 7798 5951 8114 5952
rect 11500 6016 11816 6017
rect 11500 5952 11506 6016
rect 11570 5952 11586 6016
rect 11650 5952 11666 6016
rect 11730 5952 11746 6016
rect 11810 5952 11816 6016
rect 11500 5951 11816 5952
rect 15202 6016 15518 6017
rect 15202 5952 15208 6016
rect 15272 5952 15288 6016
rect 15352 5952 15368 6016
rect 15432 5952 15448 6016
rect 15512 5952 15518 6016
rect 15202 5951 15518 5952
rect 15600 5813 16000 5840
rect 8385 5810 8451 5813
rect 11881 5810 11947 5813
rect 13905 5810 13971 5813
rect 8385 5808 13971 5810
rect 8385 5752 8390 5808
rect 8446 5752 11886 5808
rect 11942 5752 13910 5808
rect 13966 5752 13971 5808
rect 8385 5750 13971 5752
rect 8385 5747 8451 5750
rect 11881 5747 11947 5750
rect 13905 5747 13971 5750
rect 15561 5808 16000 5813
rect 15561 5752 15566 5808
rect 15622 5752 16000 5808
rect 15561 5747 16000 5752
rect 15600 5720 16000 5747
rect 2245 5472 2561 5473
rect 2245 5408 2251 5472
rect 2315 5408 2331 5472
rect 2395 5408 2411 5472
rect 2475 5408 2491 5472
rect 2555 5408 2561 5472
rect 2245 5407 2561 5408
rect 5947 5472 6263 5473
rect 5947 5408 5953 5472
rect 6017 5408 6033 5472
rect 6097 5408 6113 5472
rect 6177 5408 6193 5472
rect 6257 5408 6263 5472
rect 5947 5407 6263 5408
rect 9649 5472 9965 5473
rect 9649 5408 9655 5472
rect 9719 5408 9735 5472
rect 9799 5408 9815 5472
rect 9879 5408 9895 5472
rect 9959 5408 9965 5472
rect 9649 5407 9965 5408
rect 13351 5472 13667 5473
rect 13351 5408 13357 5472
rect 13421 5408 13437 5472
rect 13501 5408 13517 5472
rect 13581 5408 13597 5472
rect 13661 5408 13667 5472
rect 13351 5407 13667 5408
rect 15600 4992 16000 5024
rect 15600 4936 15934 4992
rect 15990 4936 16000 4992
rect 4096 4928 4412 4929
rect 4096 4864 4102 4928
rect 4166 4864 4182 4928
rect 4246 4864 4262 4928
rect 4326 4864 4342 4928
rect 4406 4864 4412 4928
rect 4096 4863 4412 4864
rect 7798 4928 8114 4929
rect 7798 4864 7804 4928
rect 7868 4864 7884 4928
rect 7948 4864 7964 4928
rect 8028 4864 8044 4928
rect 8108 4864 8114 4928
rect 7798 4863 8114 4864
rect 11500 4928 11816 4929
rect 11500 4864 11506 4928
rect 11570 4864 11586 4928
rect 11650 4864 11666 4928
rect 11730 4864 11746 4928
rect 11810 4864 11816 4928
rect 11500 4863 11816 4864
rect 15202 4928 15518 4929
rect 15202 4864 15208 4928
rect 15272 4864 15288 4928
rect 15352 4864 15368 4928
rect 15432 4864 15448 4928
rect 15512 4864 15518 4928
rect 15600 4904 16000 4936
rect 15202 4863 15518 4864
rect 2245 4384 2561 4385
rect 2245 4320 2251 4384
rect 2315 4320 2331 4384
rect 2395 4320 2411 4384
rect 2475 4320 2491 4384
rect 2555 4320 2561 4384
rect 2245 4319 2561 4320
rect 5947 4384 6263 4385
rect 5947 4320 5953 4384
rect 6017 4320 6033 4384
rect 6097 4320 6113 4384
rect 6177 4320 6193 4384
rect 6257 4320 6263 4384
rect 5947 4319 6263 4320
rect 9649 4384 9965 4385
rect 9649 4320 9655 4384
rect 9719 4320 9735 4384
rect 9799 4320 9815 4384
rect 9879 4320 9895 4384
rect 9959 4320 9965 4384
rect 9649 4319 9965 4320
rect 13351 4384 13667 4385
rect 13351 4320 13357 4384
rect 13421 4320 13437 4384
rect 13501 4320 13517 4384
rect 13581 4320 13597 4384
rect 13661 4320 13667 4384
rect 13351 4319 13667 4320
rect 13077 4178 13143 4181
rect 13905 4178 13971 4181
rect 13077 4176 13971 4178
rect 13077 4120 13082 4176
rect 13138 4120 13910 4176
rect 13966 4120 13971 4176
rect 13077 4118 13971 4120
rect 13077 4115 13143 4118
rect 13905 4115 13971 4118
rect 15009 4178 15075 4181
rect 15600 4178 16000 4208
rect 15009 4176 16000 4178
rect 15009 4120 15014 4176
rect 15070 4120 16000 4176
rect 15009 4118 16000 4120
rect 15009 4115 15075 4118
rect 15600 4088 16000 4118
rect 4096 3840 4412 3841
rect 4096 3776 4102 3840
rect 4166 3776 4182 3840
rect 4246 3776 4262 3840
rect 4326 3776 4342 3840
rect 4406 3776 4412 3840
rect 4096 3775 4412 3776
rect 7798 3840 8114 3841
rect 7798 3776 7804 3840
rect 7868 3776 7884 3840
rect 7948 3776 7964 3840
rect 8028 3776 8044 3840
rect 8108 3776 8114 3840
rect 7798 3775 8114 3776
rect 11500 3840 11816 3841
rect 11500 3776 11506 3840
rect 11570 3776 11586 3840
rect 11650 3776 11666 3840
rect 11730 3776 11746 3840
rect 11810 3776 11816 3840
rect 11500 3775 11816 3776
rect 15202 3840 15518 3841
rect 15202 3776 15208 3840
rect 15272 3776 15288 3840
rect 15352 3776 15368 3840
rect 15432 3776 15448 3840
rect 15512 3776 15518 3840
rect 15202 3775 15518 3776
rect 15009 3362 15075 3365
rect 15600 3362 16000 3392
rect 15009 3360 16000 3362
rect 15009 3304 15014 3360
rect 15070 3304 16000 3360
rect 15009 3302 16000 3304
rect 15009 3299 15075 3302
rect 2245 3296 2561 3297
rect 2245 3232 2251 3296
rect 2315 3232 2331 3296
rect 2395 3232 2411 3296
rect 2475 3232 2491 3296
rect 2555 3232 2561 3296
rect 2245 3231 2561 3232
rect 5947 3296 6263 3297
rect 5947 3232 5953 3296
rect 6017 3232 6033 3296
rect 6097 3232 6113 3296
rect 6177 3232 6193 3296
rect 6257 3232 6263 3296
rect 5947 3231 6263 3232
rect 9649 3296 9965 3297
rect 9649 3232 9655 3296
rect 9719 3232 9735 3296
rect 9799 3232 9815 3296
rect 9879 3232 9895 3296
rect 9959 3232 9965 3296
rect 9649 3231 9965 3232
rect 13351 3296 13667 3297
rect 13351 3232 13357 3296
rect 13421 3232 13437 3296
rect 13501 3232 13517 3296
rect 13581 3232 13597 3296
rect 13661 3232 13667 3296
rect 15600 3272 16000 3302
rect 13351 3231 13667 3232
rect 4096 2752 4412 2753
rect 4096 2688 4102 2752
rect 4166 2688 4182 2752
rect 4246 2688 4262 2752
rect 4326 2688 4342 2752
rect 4406 2688 4412 2752
rect 4096 2687 4412 2688
rect 7798 2752 8114 2753
rect 7798 2688 7804 2752
rect 7868 2688 7884 2752
rect 7948 2688 7964 2752
rect 8028 2688 8044 2752
rect 8108 2688 8114 2752
rect 7798 2687 8114 2688
rect 11500 2752 11816 2753
rect 11500 2688 11506 2752
rect 11570 2688 11586 2752
rect 11650 2688 11666 2752
rect 11730 2688 11746 2752
rect 11810 2688 11816 2752
rect 11500 2687 11816 2688
rect 15202 2752 15518 2753
rect 15202 2688 15208 2752
rect 15272 2688 15288 2752
rect 15352 2688 15368 2752
rect 15432 2688 15448 2752
rect 15512 2688 15518 2752
rect 15202 2687 15518 2688
rect 8293 2546 8359 2549
rect 15009 2546 15075 2549
rect 15600 2546 16000 2576
rect 8293 2544 16000 2546
rect 8293 2488 8298 2544
rect 8354 2488 15014 2544
rect 15070 2488 16000 2544
rect 8293 2486 16000 2488
rect 8293 2483 8359 2486
rect 15009 2483 15075 2486
rect 15600 2456 16000 2486
rect 2245 2208 2561 2209
rect 2245 2144 2251 2208
rect 2315 2144 2331 2208
rect 2395 2144 2411 2208
rect 2475 2144 2491 2208
rect 2555 2144 2561 2208
rect 2245 2143 2561 2144
rect 5947 2208 6263 2209
rect 5947 2144 5953 2208
rect 6017 2144 6033 2208
rect 6097 2144 6113 2208
rect 6177 2144 6193 2208
rect 6257 2144 6263 2208
rect 5947 2143 6263 2144
rect 9649 2208 9965 2209
rect 9649 2144 9655 2208
rect 9719 2144 9735 2208
rect 9799 2144 9815 2208
rect 9879 2144 9895 2208
rect 9959 2144 9965 2208
rect 9649 2143 9965 2144
rect 13351 2208 13667 2209
rect 13351 2144 13357 2208
rect 13421 2144 13437 2208
rect 13501 2144 13517 2208
rect 13581 2144 13597 2208
rect 13661 2144 13667 2208
rect 13351 2143 13667 2144
rect 10041 1866 10107 1869
rect 15009 1866 15075 1869
rect 10041 1864 15075 1866
rect 10041 1808 10046 1864
rect 10102 1808 15014 1864
rect 15070 1808 15075 1864
rect 10041 1806 15075 1808
rect 10041 1803 10107 1806
rect 15009 1803 15075 1806
rect 15600 1728 16000 1760
rect 15600 1672 15658 1728
rect 15714 1672 16000 1728
rect 4096 1664 4412 1665
rect 4096 1600 4102 1664
rect 4166 1600 4182 1664
rect 4246 1600 4262 1664
rect 4326 1600 4342 1664
rect 4406 1600 4412 1664
rect 4096 1599 4412 1600
rect 7798 1664 8114 1665
rect 7798 1600 7804 1664
rect 7868 1600 7884 1664
rect 7948 1600 7964 1664
rect 8028 1600 8044 1664
rect 8108 1600 8114 1664
rect 7798 1599 8114 1600
rect 11500 1664 11816 1665
rect 11500 1600 11506 1664
rect 11570 1600 11586 1664
rect 11650 1600 11666 1664
rect 11730 1600 11746 1664
rect 11810 1600 11816 1664
rect 11500 1599 11816 1600
rect 15202 1664 15518 1665
rect 15202 1600 15208 1664
rect 15272 1600 15288 1664
rect 15352 1600 15368 1664
rect 15432 1600 15448 1664
rect 15512 1600 15518 1664
rect 15600 1640 16000 1672
rect 15202 1599 15518 1600
rect 2245 1120 2561 1121
rect 2245 1056 2251 1120
rect 2315 1056 2331 1120
rect 2395 1056 2411 1120
rect 2475 1056 2491 1120
rect 2555 1056 2561 1120
rect 2245 1055 2561 1056
rect 5947 1120 6263 1121
rect 5947 1056 5953 1120
rect 6017 1056 6033 1120
rect 6097 1056 6113 1120
rect 6177 1056 6193 1120
rect 6257 1056 6263 1120
rect 5947 1055 6263 1056
rect 9649 1120 9965 1121
rect 9649 1056 9655 1120
rect 9719 1056 9735 1120
rect 9799 1056 9815 1120
rect 9879 1056 9895 1120
rect 9959 1056 9965 1120
rect 9649 1055 9965 1056
rect 13351 1120 13667 1121
rect 13351 1056 13357 1120
rect 13421 1056 13437 1120
rect 13501 1056 13517 1120
rect 13581 1056 13597 1120
rect 13661 1056 13667 1120
rect 13351 1055 13667 1056
rect 4096 576 4412 577
rect 4096 512 4102 576
rect 4166 512 4182 576
rect 4246 512 4262 576
rect 4326 512 4342 576
rect 4406 512 4412 576
rect 4096 511 4412 512
rect 7798 576 8114 577
rect 7798 512 7804 576
rect 7868 512 7884 576
rect 7948 512 7964 576
rect 8028 512 8044 576
rect 8108 512 8114 576
rect 7798 511 8114 512
rect 11500 576 11816 577
rect 11500 512 11506 576
rect 11570 512 11586 576
rect 11650 512 11666 576
rect 11730 512 11746 576
rect 11810 512 11816 576
rect 11500 511 11816 512
rect 15202 576 15518 577
rect 15202 512 15208 576
rect 15272 512 15288 576
rect 15352 512 15368 576
rect 15432 512 15448 576
rect 15512 512 15518 576
rect 15202 511 15518 512
<< via3 >>
rect 2251 15260 2315 15264
rect 2251 15204 2255 15260
rect 2255 15204 2311 15260
rect 2311 15204 2315 15260
rect 2251 15200 2315 15204
rect 2331 15260 2395 15264
rect 2331 15204 2335 15260
rect 2335 15204 2391 15260
rect 2391 15204 2395 15260
rect 2331 15200 2395 15204
rect 2411 15260 2475 15264
rect 2411 15204 2415 15260
rect 2415 15204 2471 15260
rect 2471 15204 2475 15260
rect 2411 15200 2475 15204
rect 2491 15260 2555 15264
rect 2491 15204 2495 15260
rect 2495 15204 2551 15260
rect 2551 15204 2555 15260
rect 2491 15200 2555 15204
rect 5953 15260 6017 15264
rect 5953 15204 5957 15260
rect 5957 15204 6013 15260
rect 6013 15204 6017 15260
rect 5953 15200 6017 15204
rect 6033 15260 6097 15264
rect 6033 15204 6037 15260
rect 6037 15204 6093 15260
rect 6093 15204 6097 15260
rect 6033 15200 6097 15204
rect 6113 15260 6177 15264
rect 6113 15204 6117 15260
rect 6117 15204 6173 15260
rect 6173 15204 6177 15260
rect 6113 15200 6177 15204
rect 6193 15260 6257 15264
rect 6193 15204 6197 15260
rect 6197 15204 6253 15260
rect 6253 15204 6257 15260
rect 6193 15200 6257 15204
rect 9655 15260 9719 15264
rect 9655 15204 9659 15260
rect 9659 15204 9715 15260
rect 9715 15204 9719 15260
rect 9655 15200 9719 15204
rect 9735 15260 9799 15264
rect 9735 15204 9739 15260
rect 9739 15204 9795 15260
rect 9795 15204 9799 15260
rect 9735 15200 9799 15204
rect 9815 15260 9879 15264
rect 9815 15204 9819 15260
rect 9819 15204 9875 15260
rect 9875 15204 9879 15260
rect 9815 15200 9879 15204
rect 9895 15260 9959 15264
rect 9895 15204 9899 15260
rect 9899 15204 9955 15260
rect 9955 15204 9959 15260
rect 9895 15200 9959 15204
rect 13357 15260 13421 15264
rect 13357 15204 13361 15260
rect 13361 15204 13417 15260
rect 13417 15204 13421 15260
rect 13357 15200 13421 15204
rect 13437 15260 13501 15264
rect 13437 15204 13441 15260
rect 13441 15204 13497 15260
rect 13497 15204 13501 15260
rect 13437 15200 13501 15204
rect 13517 15260 13581 15264
rect 13517 15204 13521 15260
rect 13521 15204 13577 15260
rect 13577 15204 13581 15260
rect 13517 15200 13581 15204
rect 13597 15260 13661 15264
rect 13597 15204 13601 15260
rect 13601 15204 13657 15260
rect 13657 15204 13661 15260
rect 13597 15200 13661 15204
rect 4102 14716 4166 14720
rect 4102 14660 4106 14716
rect 4106 14660 4162 14716
rect 4162 14660 4166 14716
rect 4102 14656 4166 14660
rect 4182 14716 4246 14720
rect 4182 14660 4186 14716
rect 4186 14660 4242 14716
rect 4242 14660 4246 14716
rect 4182 14656 4246 14660
rect 4262 14716 4326 14720
rect 4262 14660 4266 14716
rect 4266 14660 4322 14716
rect 4322 14660 4326 14716
rect 4262 14656 4326 14660
rect 4342 14716 4406 14720
rect 4342 14660 4346 14716
rect 4346 14660 4402 14716
rect 4402 14660 4406 14716
rect 4342 14656 4406 14660
rect 7804 14716 7868 14720
rect 7804 14660 7808 14716
rect 7808 14660 7864 14716
rect 7864 14660 7868 14716
rect 7804 14656 7868 14660
rect 7884 14716 7948 14720
rect 7884 14660 7888 14716
rect 7888 14660 7944 14716
rect 7944 14660 7948 14716
rect 7884 14656 7948 14660
rect 7964 14716 8028 14720
rect 7964 14660 7968 14716
rect 7968 14660 8024 14716
rect 8024 14660 8028 14716
rect 7964 14656 8028 14660
rect 8044 14716 8108 14720
rect 8044 14660 8048 14716
rect 8048 14660 8104 14716
rect 8104 14660 8108 14716
rect 8044 14656 8108 14660
rect 11506 14716 11570 14720
rect 11506 14660 11510 14716
rect 11510 14660 11566 14716
rect 11566 14660 11570 14716
rect 11506 14656 11570 14660
rect 11586 14716 11650 14720
rect 11586 14660 11590 14716
rect 11590 14660 11646 14716
rect 11646 14660 11650 14716
rect 11586 14656 11650 14660
rect 11666 14716 11730 14720
rect 11666 14660 11670 14716
rect 11670 14660 11726 14716
rect 11726 14660 11730 14716
rect 11666 14656 11730 14660
rect 11746 14716 11810 14720
rect 11746 14660 11750 14716
rect 11750 14660 11806 14716
rect 11806 14660 11810 14716
rect 11746 14656 11810 14660
rect 15208 14716 15272 14720
rect 15208 14660 15212 14716
rect 15212 14660 15268 14716
rect 15268 14660 15272 14716
rect 15208 14656 15272 14660
rect 15288 14716 15352 14720
rect 15288 14660 15292 14716
rect 15292 14660 15348 14716
rect 15348 14660 15352 14716
rect 15288 14656 15352 14660
rect 15368 14716 15432 14720
rect 15368 14660 15372 14716
rect 15372 14660 15428 14716
rect 15428 14660 15432 14716
rect 15368 14656 15432 14660
rect 15448 14716 15512 14720
rect 15448 14660 15452 14716
rect 15452 14660 15508 14716
rect 15508 14660 15512 14716
rect 15448 14656 15512 14660
rect 2251 14172 2315 14176
rect 2251 14116 2255 14172
rect 2255 14116 2311 14172
rect 2311 14116 2315 14172
rect 2251 14112 2315 14116
rect 2331 14172 2395 14176
rect 2331 14116 2335 14172
rect 2335 14116 2391 14172
rect 2391 14116 2395 14172
rect 2331 14112 2395 14116
rect 2411 14172 2475 14176
rect 2411 14116 2415 14172
rect 2415 14116 2471 14172
rect 2471 14116 2475 14172
rect 2411 14112 2475 14116
rect 2491 14172 2555 14176
rect 2491 14116 2495 14172
rect 2495 14116 2551 14172
rect 2551 14116 2555 14172
rect 2491 14112 2555 14116
rect 5953 14172 6017 14176
rect 5953 14116 5957 14172
rect 5957 14116 6013 14172
rect 6013 14116 6017 14172
rect 5953 14112 6017 14116
rect 6033 14172 6097 14176
rect 6033 14116 6037 14172
rect 6037 14116 6093 14172
rect 6093 14116 6097 14172
rect 6033 14112 6097 14116
rect 6113 14172 6177 14176
rect 6113 14116 6117 14172
rect 6117 14116 6173 14172
rect 6173 14116 6177 14172
rect 6113 14112 6177 14116
rect 6193 14172 6257 14176
rect 6193 14116 6197 14172
rect 6197 14116 6253 14172
rect 6253 14116 6257 14172
rect 6193 14112 6257 14116
rect 9655 14172 9719 14176
rect 9655 14116 9659 14172
rect 9659 14116 9715 14172
rect 9715 14116 9719 14172
rect 9655 14112 9719 14116
rect 9735 14172 9799 14176
rect 9735 14116 9739 14172
rect 9739 14116 9795 14172
rect 9795 14116 9799 14172
rect 9735 14112 9799 14116
rect 9815 14172 9879 14176
rect 9815 14116 9819 14172
rect 9819 14116 9875 14172
rect 9875 14116 9879 14172
rect 9815 14112 9879 14116
rect 9895 14172 9959 14176
rect 9895 14116 9899 14172
rect 9899 14116 9955 14172
rect 9955 14116 9959 14172
rect 9895 14112 9959 14116
rect 13357 14172 13421 14176
rect 13357 14116 13361 14172
rect 13361 14116 13417 14172
rect 13417 14116 13421 14172
rect 13357 14112 13421 14116
rect 13437 14172 13501 14176
rect 13437 14116 13441 14172
rect 13441 14116 13497 14172
rect 13497 14116 13501 14172
rect 13437 14112 13501 14116
rect 13517 14172 13581 14176
rect 13517 14116 13521 14172
rect 13521 14116 13577 14172
rect 13577 14116 13581 14172
rect 13517 14112 13581 14116
rect 13597 14172 13661 14176
rect 13597 14116 13601 14172
rect 13601 14116 13657 14172
rect 13657 14116 13661 14172
rect 13597 14112 13661 14116
rect 4102 13628 4166 13632
rect 4102 13572 4106 13628
rect 4106 13572 4162 13628
rect 4162 13572 4166 13628
rect 4102 13568 4166 13572
rect 4182 13628 4246 13632
rect 4182 13572 4186 13628
rect 4186 13572 4242 13628
rect 4242 13572 4246 13628
rect 4182 13568 4246 13572
rect 4262 13628 4326 13632
rect 4262 13572 4266 13628
rect 4266 13572 4322 13628
rect 4322 13572 4326 13628
rect 4262 13568 4326 13572
rect 4342 13628 4406 13632
rect 4342 13572 4346 13628
rect 4346 13572 4402 13628
rect 4402 13572 4406 13628
rect 4342 13568 4406 13572
rect 7804 13628 7868 13632
rect 7804 13572 7808 13628
rect 7808 13572 7864 13628
rect 7864 13572 7868 13628
rect 7804 13568 7868 13572
rect 7884 13628 7948 13632
rect 7884 13572 7888 13628
rect 7888 13572 7944 13628
rect 7944 13572 7948 13628
rect 7884 13568 7948 13572
rect 7964 13628 8028 13632
rect 7964 13572 7968 13628
rect 7968 13572 8024 13628
rect 8024 13572 8028 13628
rect 7964 13568 8028 13572
rect 8044 13628 8108 13632
rect 8044 13572 8048 13628
rect 8048 13572 8104 13628
rect 8104 13572 8108 13628
rect 8044 13568 8108 13572
rect 11506 13628 11570 13632
rect 11506 13572 11510 13628
rect 11510 13572 11566 13628
rect 11566 13572 11570 13628
rect 11506 13568 11570 13572
rect 11586 13628 11650 13632
rect 11586 13572 11590 13628
rect 11590 13572 11646 13628
rect 11646 13572 11650 13628
rect 11586 13568 11650 13572
rect 11666 13628 11730 13632
rect 11666 13572 11670 13628
rect 11670 13572 11726 13628
rect 11726 13572 11730 13628
rect 11666 13568 11730 13572
rect 11746 13628 11810 13632
rect 11746 13572 11750 13628
rect 11750 13572 11806 13628
rect 11806 13572 11810 13628
rect 11746 13568 11810 13572
rect 15208 13628 15272 13632
rect 15208 13572 15212 13628
rect 15212 13572 15268 13628
rect 15268 13572 15272 13628
rect 15208 13568 15272 13572
rect 15288 13628 15352 13632
rect 15288 13572 15292 13628
rect 15292 13572 15348 13628
rect 15348 13572 15352 13628
rect 15288 13568 15352 13572
rect 15368 13628 15432 13632
rect 15368 13572 15372 13628
rect 15372 13572 15428 13628
rect 15428 13572 15432 13628
rect 15368 13568 15432 13572
rect 15448 13628 15512 13632
rect 15448 13572 15452 13628
rect 15452 13572 15508 13628
rect 15508 13572 15512 13628
rect 15448 13568 15512 13572
rect 2251 13084 2315 13088
rect 2251 13028 2255 13084
rect 2255 13028 2311 13084
rect 2311 13028 2315 13084
rect 2251 13024 2315 13028
rect 2331 13084 2395 13088
rect 2331 13028 2335 13084
rect 2335 13028 2391 13084
rect 2391 13028 2395 13084
rect 2331 13024 2395 13028
rect 2411 13084 2475 13088
rect 2411 13028 2415 13084
rect 2415 13028 2471 13084
rect 2471 13028 2475 13084
rect 2411 13024 2475 13028
rect 2491 13084 2555 13088
rect 2491 13028 2495 13084
rect 2495 13028 2551 13084
rect 2551 13028 2555 13084
rect 2491 13024 2555 13028
rect 5953 13084 6017 13088
rect 5953 13028 5957 13084
rect 5957 13028 6013 13084
rect 6013 13028 6017 13084
rect 5953 13024 6017 13028
rect 6033 13084 6097 13088
rect 6033 13028 6037 13084
rect 6037 13028 6093 13084
rect 6093 13028 6097 13084
rect 6033 13024 6097 13028
rect 6113 13084 6177 13088
rect 6113 13028 6117 13084
rect 6117 13028 6173 13084
rect 6173 13028 6177 13084
rect 6113 13024 6177 13028
rect 6193 13084 6257 13088
rect 6193 13028 6197 13084
rect 6197 13028 6253 13084
rect 6253 13028 6257 13084
rect 6193 13024 6257 13028
rect 9655 13084 9719 13088
rect 9655 13028 9659 13084
rect 9659 13028 9715 13084
rect 9715 13028 9719 13084
rect 9655 13024 9719 13028
rect 9735 13084 9799 13088
rect 9735 13028 9739 13084
rect 9739 13028 9795 13084
rect 9795 13028 9799 13084
rect 9735 13024 9799 13028
rect 9815 13084 9879 13088
rect 9815 13028 9819 13084
rect 9819 13028 9875 13084
rect 9875 13028 9879 13084
rect 9815 13024 9879 13028
rect 9895 13084 9959 13088
rect 9895 13028 9899 13084
rect 9899 13028 9955 13084
rect 9955 13028 9959 13084
rect 9895 13024 9959 13028
rect 13357 13084 13421 13088
rect 13357 13028 13361 13084
rect 13361 13028 13417 13084
rect 13417 13028 13421 13084
rect 13357 13024 13421 13028
rect 13437 13084 13501 13088
rect 13437 13028 13441 13084
rect 13441 13028 13497 13084
rect 13497 13028 13501 13084
rect 13437 13024 13501 13028
rect 13517 13084 13581 13088
rect 13517 13028 13521 13084
rect 13521 13028 13577 13084
rect 13577 13028 13581 13084
rect 13517 13024 13581 13028
rect 13597 13084 13661 13088
rect 13597 13028 13601 13084
rect 13601 13028 13657 13084
rect 13657 13028 13661 13084
rect 13597 13024 13661 13028
rect 4102 12540 4166 12544
rect 4102 12484 4106 12540
rect 4106 12484 4162 12540
rect 4162 12484 4166 12540
rect 4102 12480 4166 12484
rect 4182 12540 4246 12544
rect 4182 12484 4186 12540
rect 4186 12484 4242 12540
rect 4242 12484 4246 12540
rect 4182 12480 4246 12484
rect 4262 12540 4326 12544
rect 4262 12484 4266 12540
rect 4266 12484 4322 12540
rect 4322 12484 4326 12540
rect 4262 12480 4326 12484
rect 4342 12540 4406 12544
rect 4342 12484 4346 12540
rect 4346 12484 4402 12540
rect 4402 12484 4406 12540
rect 4342 12480 4406 12484
rect 7804 12540 7868 12544
rect 7804 12484 7808 12540
rect 7808 12484 7864 12540
rect 7864 12484 7868 12540
rect 7804 12480 7868 12484
rect 7884 12540 7948 12544
rect 7884 12484 7888 12540
rect 7888 12484 7944 12540
rect 7944 12484 7948 12540
rect 7884 12480 7948 12484
rect 7964 12540 8028 12544
rect 7964 12484 7968 12540
rect 7968 12484 8024 12540
rect 8024 12484 8028 12540
rect 7964 12480 8028 12484
rect 8044 12540 8108 12544
rect 8044 12484 8048 12540
rect 8048 12484 8104 12540
rect 8104 12484 8108 12540
rect 8044 12480 8108 12484
rect 11506 12540 11570 12544
rect 11506 12484 11510 12540
rect 11510 12484 11566 12540
rect 11566 12484 11570 12540
rect 11506 12480 11570 12484
rect 11586 12540 11650 12544
rect 11586 12484 11590 12540
rect 11590 12484 11646 12540
rect 11646 12484 11650 12540
rect 11586 12480 11650 12484
rect 11666 12540 11730 12544
rect 11666 12484 11670 12540
rect 11670 12484 11726 12540
rect 11726 12484 11730 12540
rect 11666 12480 11730 12484
rect 11746 12540 11810 12544
rect 11746 12484 11750 12540
rect 11750 12484 11806 12540
rect 11806 12484 11810 12540
rect 11746 12480 11810 12484
rect 15208 12540 15272 12544
rect 15208 12484 15212 12540
rect 15212 12484 15268 12540
rect 15268 12484 15272 12540
rect 15208 12480 15272 12484
rect 15288 12540 15352 12544
rect 15288 12484 15292 12540
rect 15292 12484 15348 12540
rect 15348 12484 15352 12540
rect 15288 12480 15352 12484
rect 15368 12540 15432 12544
rect 15368 12484 15372 12540
rect 15372 12484 15428 12540
rect 15428 12484 15432 12540
rect 15368 12480 15432 12484
rect 15448 12540 15512 12544
rect 15448 12484 15452 12540
rect 15452 12484 15508 12540
rect 15508 12484 15512 12540
rect 15448 12480 15512 12484
rect 2251 11996 2315 12000
rect 2251 11940 2255 11996
rect 2255 11940 2311 11996
rect 2311 11940 2315 11996
rect 2251 11936 2315 11940
rect 2331 11996 2395 12000
rect 2331 11940 2335 11996
rect 2335 11940 2391 11996
rect 2391 11940 2395 11996
rect 2331 11936 2395 11940
rect 2411 11996 2475 12000
rect 2411 11940 2415 11996
rect 2415 11940 2471 11996
rect 2471 11940 2475 11996
rect 2411 11936 2475 11940
rect 2491 11996 2555 12000
rect 2491 11940 2495 11996
rect 2495 11940 2551 11996
rect 2551 11940 2555 11996
rect 2491 11936 2555 11940
rect 5953 11996 6017 12000
rect 5953 11940 5957 11996
rect 5957 11940 6013 11996
rect 6013 11940 6017 11996
rect 5953 11936 6017 11940
rect 6033 11996 6097 12000
rect 6033 11940 6037 11996
rect 6037 11940 6093 11996
rect 6093 11940 6097 11996
rect 6033 11936 6097 11940
rect 6113 11996 6177 12000
rect 6113 11940 6117 11996
rect 6117 11940 6173 11996
rect 6173 11940 6177 11996
rect 6113 11936 6177 11940
rect 6193 11996 6257 12000
rect 6193 11940 6197 11996
rect 6197 11940 6253 11996
rect 6253 11940 6257 11996
rect 6193 11936 6257 11940
rect 9655 11996 9719 12000
rect 9655 11940 9659 11996
rect 9659 11940 9715 11996
rect 9715 11940 9719 11996
rect 9655 11936 9719 11940
rect 9735 11996 9799 12000
rect 9735 11940 9739 11996
rect 9739 11940 9795 11996
rect 9795 11940 9799 11996
rect 9735 11936 9799 11940
rect 9815 11996 9879 12000
rect 9815 11940 9819 11996
rect 9819 11940 9875 11996
rect 9875 11940 9879 11996
rect 9815 11936 9879 11940
rect 9895 11996 9959 12000
rect 9895 11940 9899 11996
rect 9899 11940 9955 11996
rect 9955 11940 9959 11996
rect 9895 11936 9959 11940
rect 13357 11996 13421 12000
rect 13357 11940 13361 11996
rect 13361 11940 13417 11996
rect 13417 11940 13421 11996
rect 13357 11936 13421 11940
rect 13437 11996 13501 12000
rect 13437 11940 13441 11996
rect 13441 11940 13497 11996
rect 13497 11940 13501 11996
rect 13437 11936 13501 11940
rect 13517 11996 13581 12000
rect 13517 11940 13521 11996
rect 13521 11940 13577 11996
rect 13577 11940 13581 11996
rect 13517 11936 13581 11940
rect 13597 11996 13661 12000
rect 13597 11940 13601 11996
rect 13601 11940 13657 11996
rect 13657 11940 13661 11996
rect 13597 11936 13661 11940
rect 4102 11452 4166 11456
rect 4102 11396 4106 11452
rect 4106 11396 4162 11452
rect 4162 11396 4166 11452
rect 4102 11392 4166 11396
rect 4182 11452 4246 11456
rect 4182 11396 4186 11452
rect 4186 11396 4242 11452
rect 4242 11396 4246 11452
rect 4182 11392 4246 11396
rect 4262 11452 4326 11456
rect 4262 11396 4266 11452
rect 4266 11396 4322 11452
rect 4322 11396 4326 11452
rect 4262 11392 4326 11396
rect 4342 11452 4406 11456
rect 4342 11396 4346 11452
rect 4346 11396 4402 11452
rect 4402 11396 4406 11452
rect 4342 11392 4406 11396
rect 7804 11452 7868 11456
rect 7804 11396 7808 11452
rect 7808 11396 7864 11452
rect 7864 11396 7868 11452
rect 7804 11392 7868 11396
rect 7884 11452 7948 11456
rect 7884 11396 7888 11452
rect 7888 11396 7944 11452
rect 7944 11396 7948 11452
rect 7884 11392 7948 11396
rect 7964 11452 8028 11456
rect 7964 11396 7968 11452
rect 7968 11396 8024 11452
rect 8024 11396 8028 11452
rect 7964 11392 8028 11396
rect 8044 11452 8108 11456
rect 8044 11396 8048 11452
rect 8048 11396 8104 11452
rect 8104 11396 8108 11452
rect 8044 11392 8108 11396
rect 11506 11452 11570 11456
rect 11506 11396 11510 11452
rect 11510 11396 11566 11452
rect 11566 11396 11570 11452
rect 11506 11392 11570 11396
rect 11586 11452 11650 11456
rect 11586 11396 11590 11452
rect 11590 11396 11646 11452
rect 11646 11396 11650 11452
rect 11586 11392 11650 11396
rect 11666 11452 11730 11456
rect 11666 11396 11670 11452
rect 11670 11396 11726 11452
rect 11726 11396 11730 11452
rect 11666 11392 11730 11396
rect 11746 11452 11810 11456
rect 11746 11396 11750 11452
rect 11750 11396 11806 11452
rect 11806 11396 11810 11452
rect 11746 11392 11810 11396
rect 15208 11452 15272 11456
rect 15208 11396 15212 11452
rect 15212 11396 15268 11452
rect 15268 11396 15272 11452
rect 15208 11392 15272 11396
rect 15288 11452 15352 11456
rect 15288 11396 15292 11452
rect 15292 11396 15348 11452
rect 15348 11396 15352 11452
rect 15288 11392 15352 11396
rect 15368 11452 15432 11456
rect 15368 11396 15372 11452
rect 15372 11396 15428 11452
rect 15428 11396 15432 11452
rect 15368 11392 15432 11396
rect 15448 11452 15512 11456
rect 15448 11396 15452 11452
rect 15452 11396 15508 11452
rect 15508 11396 15512 11452
rect 15448 11392 15512 11396
rect 2251 10908 2315 10912
rect 2251 10852 2255 10908
rect 2255 10852 2311 10908
rect 2311 10852 2315 10908
rect 2251 10848 2315 10852
rect 2331 10908 2395 10912
rect 2331 10852 2335 10908
rect 2335 10852 2391 10908
rect 2391 10852 2395 10908
rect 2331 10848 2395 10852
rect 2411 10908 2475 10912
rect 2411 10852 2415 10908
rect 2415 10852 2471 10908
rect 2471 10852 2475 10908
rect 2411 10848 2475 10852
rect 2491 10908 2555 10912
rect 2491 10852 2495 10908
rect 2495 10852 2551 10908
rect 2551 10852 2555 10908
rect 2491 10848 2555 10852
rect 5953 10908 6017 10912
rect 5953 10852 5957 10908
rect 5957 10852 6013 10908
rect 6013 10852 6017 10908
rect 5953 10848 6017 10852
rect 6033 10908 6097 10912
rect 6033 10852 6037 10908
rect 6037 10852 6093 10908
rect 6093 10852 6097 10908
rect 6033 10848 6097 10852
rect 6113 10908 6177 10912
rect 6113 10852 6117 10908
rect 6117 10852 6173 10908
rect 6173 10852 6177 10908
rect 6113 10848 6177 10852
rect 6193 10908 6257 10912
rect 6193 10852 6197 10908
rect 6197 10852 6253 10908
rect 6253 10852 6257 10908
rect 6193 10848 6257 10852
rect 9655 10908 9719 10912
rect 9655 10852 9659 10908
rect 9659 10852 9715 10908
rect 9715 10852 9719 10908
rect 9655 10848 9719 10852
rect 9735 10908 9799 10912
rect 9735 10852 9739 10908
rect 9739 10852 9795 10908
rect 9795 10852 9799 10908
rect 9735 10848 9799 10852
rect 9815 10908 9879 10912
rect 9815 10852 9819 10908
rect 9819 10852 9875 10908
rect 9875 10852 9879 10908
rect 9815 10848 9879 10852
rect 9895 10908 9959 10912
rect 9895 10852 9899 10908
rect 9899 10852 9955 10908
rect 9955 10852 9959 10908
rect 9895 10848 9959 10852
rect 13357 10908 13421 10912
rect 13357 10852 13361 10908
rect 13361 10852 13417 10908
rect 13417 10852 13421 10908
rect 13357 10848 13421 10852
rect 13437 10908 13501 10912
rect 13437 10852 13441 10908
rect 13441 10852 13497 10908
rect 13497 10852 13501 10908
rect 13437 10848 13501 10852
rect 13517 10908 13581 10912
rect 13517 10852 13521 10908
rect 13521 10852 13577 10908
rect 13577 10852 13581 10908
rect 13517 10848 13581 10852
rect 13597 10908 13661 10912
rect 13597 10852 13601 10908
rect 13601 10852 13657 10908
rect 13657 10852 13661 10908
rect 13597 10848 13661 10852
rect 4102 10364 4166 10368
rect 4102 10308 4106 10364
rect 4106 10308 4162 10364
rect 4162 10308 4166 10364
rect 4102 10304 4166 10308
rect 4182 10364 4246 10368
rect 4182 10308 4186 10364
rect 4186 10308 4242 10364
rect 4242 10308 4246 10364
rect 4182 10304 4246 10308
rect 4262 10364 4326 10368
rect 4262 10308 4266 10364
rect 4266 10308 4322 10364
rect 4322 10308 4326 10364
rect 4262 10304 4326 10308
rect 4342 10364 4406 10368
rect 4342 10308 4346 10364
rect 4346 10308 4402 10364
rect 4402 10308 4406 10364
rect 4342 10304 4406 10308
rect 7804 10364 7868 10368
rect 7804 10308 7808 10364
rect 7808 10308 7864 10364
rect 7864 10308 7868 10364
rect 7804 10304 7868 10308
rect 7884 10364 7948 10368
rect 7884 10308 7888 10364
rect 7888 10308 7944 10364
rect 7944 10308 7948 10364
rect 7884 10304 7948 10308
rect 7964 10364 8028 10368
rect 7964 10308 7968 10364
rect 7968 10308 8024 10364
rect 8024 10308 8028 10364
rect 7964 10304 8028 10308
rect 8044 10364 8108 10368
rect 8044 10308 8048 10364
rect 8048 10308 8104 10364
rect 8104 10308 8108 10364
rect 8044 10304 8108 10308
rect 11506 10364 11570 10368
rect 11506 10308 11510 10364
rect 11510 10308 11566 10364
rect 11566 10308 11570 10364
rect 11506 10304 11570 10308
rect 11586 10364 11650 10368
rect 11586 10308 11590 10364
rect 11590 10308 11646 10364
rect 11646 10308 11650 10364
rect 11586 10304 11650 10308
rect 11666 10364 11730 10368
rect 11666 10308 11670 10364
rect 11670 10308 11726 10364
rect 11726 10308 11730 10364
rect 11666 10304 11730 10308
rect 11746 10364 11810 10368
rect 11746 10308 11750 10364
rect 11750 10308 11806 10364
rect 11806 10308 11810 10364
rect 11746 10304 11810 10308
rect 15208 10364 15272 10368
rect 15208 10308 15212 10364
rect 15212 10308 15268 10364
rect 15268 10308 15272 10364
rect 15208 10304 15272 10308
rect 15288 10364 15352 10368
rect 15288 10308 15292 10364
rect 15292 10308 15348 10364
rect 15348 10308 15352 10364
rect 15288 10304 15352 10308
rect 15368 10364 15432 10368
rect 15368 10308 15372 10364
rect 15372 10308 15428 10364
rect 15428 10308 15432 10364
rect 15368 10304 15432 10308
rect 15448 10364 15512 10368
rect 15448 10308 15452 10364
rect 15452 10308 15508 10364
rect 15508 10308 15512 10364
rect 15448 10304 15512 10308
rect 2251 9820 2315 9824
rect 2251 9764 2255 9820
rect 2255 9764 2311 9820
rect 2311 9764 2315 9820
rect 2251 9760 2315 9764
rect 2331 9820 2395 9824
rect 2331 9764 2335 9820
rect 2335 9764 2391 9820
rect 2391 9764 2395 9820
rect 2331 9760 2395 9764
rect 2411 9820 2475 9824
rect 2411 9764 2415 9820
rect 2415 9764 2471 9820
rect 2471 9764 2475 9820
rect 2411 9760 2475 9764
rect 2491 9820 2555 9824
rect 2491 9764 2495 9820
rect 2495 9764 2551 9820
rect 2551 9764 2555 9820
rect 2491 9760 2555 9764
rect 5953 9820 6017 9824
rect 5953 9764 5957 9820
rect 5957 9764 6013 9820
rect 6013 9764 6017 9820
rect 5953 9760 6017 9764
rect 6033 9820 6097 9824
rect 6033 9764 6037 9820
rect 6037 9764 6093 9820
rect 6093 9764 6097 9820
rect 6033 9760 6097 9764
rect 6113 9820 6177 9824
rect 6113 9764 6117 9820
rect 6117 9764 6173 9820
rect 6173 9764 6177 9820
rect 6113 9760 6177 9764
rect 6193 9820 6257 9824
rect 6193 9764 6197 9820
rect 6197 9764 6253 9820
rect 6253 9764 6257 9820
rect 6193 9760 6257 9764
rect 9655 9820 9719 9824
rect 9655 9764 9659 9820
rect 9659 9764 9715 9820
rect 9715 9764 9719 9820
rect 9655 9760 9719 9764
rect 9735 9820 9799 9824
rect 9735 9764 9739 9820
rect 9739 9764 9795 9820
rect 9795 9764 9799 9820
rect 9735 9760 9799 9764
rect 9815 9820 9879 9824
rect 9815 9764 9819 9820
rect 9819 9764 9875 9820
rect 9875 9764 9879 9820
rect 9815 9760 9879 9764
rect 9895 9820 9959 9824
rect 9895 9764 9899 9820
rect 9899 9764 9955 9820
rect 9955 9764 9959 9820
rect 9895 9760 9959 9764
rect 13357 9820 13421 9824
rect 13357 9764 13361 9820
rect 13361 9764 13417 9820
rect 13417 9764 13421 9820
rect 13357 9760 13421 9764
rect 13437 9820 13501 9824
rect 13437 9764 13441 9820
rect 13441 9764 13497 9820
rect 13497 9764 13501 9820
rect 13437 9760 13501 9764
rect 13517 9820 13581 9824
rect 13517 9764 13521 9820
rect 13521 9764 13577 9820
rect 13577 9764 13581 9820
rect 13517 9760 13581 9764
rect 13597 9820 13661 9824
rect 13597 9764 13601 9820
rect 13601 9764 13657 9820
rect 13657 9764 13661 9820
rect 13597 9760 13661 9764
rect 4102 9276 4166 9280
rect 4102 9220 4106 9276
rect 4106 9220 4162 9276
rect 4162 9220 4166 9276
rect 4102 9216 4166 9220
rect 4182 9276 4246 9280
rect 4182 9220 4186 9276
rect 4186 9220 4242 9276
rect 4242 9220 4246 9276
rect 4182 9216 4246 9220
rect 4262 9276 4326 9280
rect 4262 9220 4266 9276
rect 4266 9220 4322 9276
rect 4322 9220 4326 9276
rect 4262 9216 4326 9220
rect 4342 9276 4406 9280
rect 4342 9220 4346 9276
rect 4346 9220 4402 9276
rect 4402 9220 4406 9276
rect 4342 9216 4406 9220
rect 7804 9276 7868 9280
rect 7804 9220 7808 9276
rect 7808 9220 7864 9276
rect 7864 9220 7868 9276
rect 7804 9216 7868 9220
rect 7884 9276 7948 9280
rect 7884 9220 7888 9276
rect 7888 9220 7944 9276
rect 7944 9220 7948 9276
rect 7884 9216 7948 9220
rect 7964 9276 8028 9280
rect 7964 9220 7968 9276
rect 7968 9220 8024 9276
rect 8024 9220 8028 9276
rect 7964 9216 8028 9220
rect 8044 9276 8108 9280
rect 8044 9220 8048 9276
rect 8048 9220 8104 9276
rect 8104 9220 8108 9276
rect 8044 9216 8108 9220
rect 11506 9276 11570 9280
rect 11506 9220 11510 9276
rect 11510 9220 11566 9276
rect 11566 9220 11570 9276
rect 11506 9216 11570 9220
rect 11586 9276 11650 9280
rect 11586 9220 11590 9276
rect 11590 9220 11646 9276
rect 11646 9220 11650 9276
rect 11586 9216 11650 9220
rect 11666 9276 11730 9280
rect 11666 9220 11670 9276
rect 11670 9220 11726 9276
rect 11726 9220 11730 9276
rect 11666 9216 11730 9220
rect 11746 9276 11810 9280
rect 11746 9220 11750 9276
rect 11750 9220 11806 9276
rect 11806 9220 11810 9276
rect 11746 9216 11810 9220
rect 15208 9276 15272 9280
rect 15208 9220 15212 9276
rect 15212 9220 15268 9276
rect 15268 9220 15272 9276
rect 15208 9216 15272 9220
rect 15288 9276 15352 9280
rect 15288 9220 15292 9276
rect 15292 9220 15348 9276
rect 15348 9220 15352 9276
rect 15288 9216 15352 9220
rect 15368 9276 15432 9280
rect 15368 9220 15372 9276
rect 15372 9220 15428 9276
rect 15428 9220 15432 9276
rect 15368 9216 15432 9220
rect 15448 9276 15512 9280
rect 15448 9220 15452 9276
rect 15452 9220 15508 9276
rect 15508 9220 15512 9276
rect 15448 9216 15512 9220
rect 2251 8732 2315 8736
rect 2251 8676 2255 8732
rect 2255 8676 2311 8732
rect 2311 8676 2315 8732
rect 2251 8672 2315 8676
rect 2331 8732 2395 8736
rect 2331 8676 2335 8732
rect 2335 8676 2391 8732
rect 2391 8676 2395 8732
rect 2331 8672 2395 8676
rect 2411 8732 2475 8736
rect 2411 8676 2415 8732
rect 2415 8676 2471 8732
rect 2471 8676 2475 8732
rect 2411 8672 2475 8676
rect 2491 8732 2555 8736
rect 2491 8676 2495 8732
rect 2495 8676 2551 8732
rect 2551 8676 2555 8732
rect 2491 8672 2555 8676
rect 5953 8732 6017 8736
rect 5953 8676 5957 8732
rect 5957 8676 6013 8732
rect 6013 8676 6017 8732
rect 5953 8672 6017 8676
rect 6033 8732 6097 8736
rect 6033 8676 6037 8732
rect 6037 8676 6093 8732
rect 6093 8676 6097 8732
rect 6033 8672 6097 8676
rect 6113 8732 6177 8736
rect 6113 8676 6117 8732
rect 6117 8676 6173 8732
rect 6173 8676 6177 8732
rect 6113 8672 6177 8676
rect 6193 8732 6257 8736
rect 6193 8676 6197 8732
rect 6197 8676 6253 8732
rect 6253 8676 6257 8732
rect 6193 8672 6257 8676
rect 9655 8732 9719 8736
rect 9655 8676 9659 8732
rect 9659 8676 9715 8732
rect 9715 8676 9719 8732
rect 9655 8672 9719 8676
rect 9735 8732 9799 8736
rect 9735 8676 9739 8732
rect 9739 8676 9795 8732
rect 9795 8676 9799 8732
rect 9735 8672 9799 8676
rect 9815 8732 9879 8736
rect 9815 8676 9819 8732
rect 9819 8676 9875 8732
rect 9875 8676 9879 8732
rect 9815 8672 9879 8676
rect 9895 8732 9959 8736
rect 9895 8676 9899 8732
rect 9899 8676 9955 8732
rect 9955 8676 9959 8732
rect 9895 8672 9959 8676
rect 13357 8732 13421 8736
rect 13357 8676 13361 8732
rect 13361 8676 13417 8732
rect 13417 8676 13421 8732
rect 13357 8672 13421 8676
rect 13437 8732 13501 8736
rect 13437 8676 13441 8732
rect 13441 8676 13497 8732
rect 13497 8676 13501 8732
rect 13437 8672 13501 8676
rect 13517 8732 13581 8736
rect 13517 8676 13521 8732
rect 13521 8676 13577 8732
rect 13577 8676 13581 8732
rect 13517 8672 13581 8676
rect 13597 8732 13661 8736
rect 13597 8676 13601 8732
rect 13601 8676 13657 8732
rect 13657 8676 13661 8732
rect 13597 8672 13661 8676
rect 4102 8188 4166 8192
rect 4102 8132 4106 8188
rect 4106 8132 4162 8188
rect 4162 8132 4166 8188
rect 4102 8128 4166 8132
rect 4182 8188 4246 8192
rect 4182 8132 4186 8188
rect 4186 8132 4242 8188
rect 4242 8132 4246 8188
rect 4182 8128 4246 8132
rect 4262 8188 4326 8192
rect 4262 8132 4266 8188
rect 4266 8132 4322 8188
rect 4322 8132 4326 8188
rect 4262 8128 4326 8132
rect 4342 8188 4406 8192
rect 4342 8132 4346 8188
rect 4346 8132 4402 8188
rect 4402 8132 4406 8188
rect 4342 8128 4406 8132
rect 7804 8188 7868 8192
rect 7804 8132 7808 8188
rect 7808 8132 7864 8188
rect 7864 8132 7868 8188
rect 7804 8128 7868 8132
rect 7884 8188 7948 8192
rect 7884 8132 7888 8188
rect 7888 8132 7944 8188
rect 7944 8132 7948 8188
rect 7884 8128 7948 8132
rect 7964 8188 8028 8192
rect 7964 8132 7968 8188
rect 7968 8132 8024 8188
rect 8024 8132 8028 8188
rect 7964 8128 8028 8132
rect 8044 8188 8108 8192
rect 8044 8132 8048 8188
rect 8048 8132 8104 8188
rect 8104 8132 8108 8188
rect 8044 8128 8108 8132
rect 11506 8188 11570 8192
rect 11506 8132 11510 8188
rect 11510 8132 11566 8188
rect 11566 8132 11570 8188
rect 11506 8128 11570 8132
rect 11586 8188 11650 8192
rect 11586 8132 11590 8188
rect 11590 8132 11646 8188
rect 11646 8132 11650 8188
rect 11586 8128 11650 8132
rect 11666 8188 11730 8192
rect 11666 8132 11670 8188
rect 11670 8132 11726 8188
rect 11726 8132 11730 8188
rect 11666 8128 11730 8132
rect 11746 8188 11810 8192
rect 11746 8132 11750 8188
rect 11750 8132 11806 8188
rect 11806 8132 11810 8188
rect 11746 8128 11810 8132
rect 15208 8188 15272 8192
rect 15208 8132 15212 8188
rect 15212 8132 15268 8188
rect 15268 8132 15272 8188
rect 15208 8128 15272 8132
rect 15288 8188 15352 8192
rect 15288 8132 15292 8188
rect 15292 8132 15348 8188
rect 15348 8132 15352 8188
rect 15288 8128 15352 8132
rect 15368 8188 15432 8192
rect 15368 8132 15372 8188
rect 15372 8132 15428 8188
rect 15428 8132 15432 8188
rect 15368 8128 15432 8132
rect 15448 8188 15512 8192
rect 15448 8132 15452 8188
rect 15452 8132 15508 8188
rect 15508 8132 15512 8188
rect 15448 8128 15512 8132
rect 2251 7644 2315 7648
rect 2251 7588 2255 7644
rect 2255 7588 2311 7644
rect 2311 7588 2315 7644
rect 2251 7584 2315 7588
rect 2331 7644 2395 7648
rect 2331 7588 2335 7644
rect 2335 7588 2391 7644
rect 2391 7588 2395 7644
rect 2331 7584 2395 7588
rect 2411 7644 2475 7648
rect 2411 7588 2415 7644
rect 2415 7588 2471 7644
rect 2471 7588 2475 7644
rect 2411 7584 2475 7588
rect 2491 7644 2555 7648
rect 2491 7588 2495 7644
rect 2495 7588 2551 7644
rect 2551 7588 2555 7644
rect 2491 7584 2555 7588
rect 5953 7644 6017 7648
rect 5953 7588 5957 7644
rect 5957 7588 6013 7644
rect 6013 7588 6017 7644
rect 5953 7584 6017 7588
rect 6033 7644 6097 7648
rect 6033 7588 6037 7644
rect 6037 7588 6093 7644
rect 6093 7588 6097 7644
rect 6033 7584 6097 7588
rect 6113 7644 6177 7648
rect 6113 7588 6117 7644
rect 6117 7588 6173 7644
rect 6173 7588 6177 7644
rect 6113 7584 6177 7588
rect 6193 7644 6257 7648
rect 6193 7588 6197 7644
rect 6197 7588 6253 7644
rect 6253 7588 6257 7644
rect 6193 7584 6257 7588
rect 9655 7644 9719 7648
rect 9655 7588 9659 7644
rect 9659 7588 9715 7644
rect 9715 7588 9719 7644
rect 9655 7584 9719 7588
rect 9735 7644 9799 7648
rect 9735 7588 9739 7644
rect 9739 7588 9795 7644
rect 9795 7588 9799 7644
rect 9735 7584 9799 7588
rect 9815 7644 9879 7648
rect 9815 7588 9819 7644
rect 9819 7588 9875 7644
rect 9875 7588 9879 7644
rect 9815 7584 9879 7588
rect 9895 7644 9959 7648
rect 9895 7588 9899 7644
rect 9899 7588 9955 7644
rect 9955 7588 9959 7644
rect 9895 7584 9959 7588
rect 13357 7644 13421 7648
rect 13357 7588 13361 7644
rect 13361 7588 13417 7644
rect 13417 7588 13421 7644
rect 13357 7584 13421 7588
rect 13437 7644 13501 7648
rect 13437 7588 13441 7644
rect 13441 7588 13497 7644
rect 13497 7588 13501 7644
rect 13437 7584 13501 7588
rect 13517 7644 13581 7648
rect 13517 7588 13521 7644
rect 13521 7588 13577 7644
rect 13577 7588 13581 7644
rect 13517 7584 13581 7588
rect 13597 7644 13661 7648
rect 13597 7588 13601 7644
rect 13601 7588 13657 7644
rect 13657 7588 13661 7644
rect 13597 7584 13661 7588
rect 4102 7100 4166 7104
rect 4102 7044 4106 7100
rect 4106 7044 4162 7100
rect 4162 7044 4166 7100
rect 4102 7040 4166 7044
rect 4182 7100 4246 7104
rect 4182 7044 4186 7100
rect 4186 7044 4242 7100
rect 4242 7044 4246 7100
rect 4182 7040 4246 7044
rect 4262 7100 4326 7104
rect 4262 7044 4266 7100
rect 4266 7044 4322 7100
rect 4322 7044 4326 7100
rect 4262 7040 4326 7044
rect 4342 7100 4406 7104
rect 4342 7044 4346 7100
rect 4346 7044 4402 7100
rect 4402 7044 4406 7100
rect 4342 7040 4406 7044
rect 7804 7100 7868 7104
rect 7804 7044 7808 7100
rect 7808 7044 7864 7100
rect 7864 7044 7868 7100
rect 7804 7040 7868 7044
rect 7884 7100 7948 7104
rect 7884 7044 7888 7100
rect 7888 7044 7944 7100
rect 7944 7044 7948 7100
rect 7884 7040 7948 7044
rect 7964 7100 8028 7104
rect 7964 7044 7968 7100
rect 7968 7044 8024 7100
rect 8024 7044 8028 7100
rect 7964 7040 8028 7044
rect 8044 7100 8108 7104
rect 8044 7044 8048 7100
rect 8048 7044 8104 7100
rect 8104 7044 8108 7100
rect 8044 7040 8108 7044
rect 11506 7100 11570 7104
rect 11506 7044 11510 7100
rect 11510 7044 11566 7100
rect 11566 7044 11570 7100
rect 11506 7040 11570 7044
rect 11586 7100 11650 7104
rect 11586 7044 11590 7100
rect 11590 7044 11646 7100
rect 11646 7044 11650 7100
rect 11586 7040 11650 7044
rect 11666 7100 11730 7104
rect 11666 7044 11670 7100
rect 11670 7044 11726 7100
rect 11726 7044 11730 7100
rect 11666 7040 11730 7044
rect 11746 7100 11810 7104
rect 11746 7044 11750 7100
rect 11750 7044 11806 7100
rect 11806 7044 11810 7100
rect 11746 7040 11810 7044
rect 15208 7100 15272 7104
rect 15208 7044 15212 7100
rect 15212 7044 15268 7100
rect 15268 7044 15272 7100
rect 15208 7040 15272 7044
rect 15288 7100 15352 7104
rect 15288 7044 15292 7100
rect 15292 7044 15348 7100
rect 15348 7044 15352 7100
rect 15288 7040 15352 7044
rect 15368 7100 15432 7104
rect 15368 7044 15372 7100
rect 15372 7044 15428 7100
rect 15428 7044 15432 7100
rect 15368 7040 15432 7044
rect 15448 7100 15512 7104
rect 15448 7044 15452 7100
rect 15452 7044 15508 7100
rect 15508 7044 15512 7100
rect 15448 7040 15512 7044
rect 2251 6556 2315 6560
rect 2251 6500 2255 6556
rect 2255 6500 2311 6556
rect 2311 6500 2315 6556
rect 2251 6496 2315 6500
rect 2331 6556 2395 6560
rect 2331 6500 2335 6556
rect 2335 6500 2391 6556
rect 2391 6500 2395 6556
rect 2331 6496 2395 6500
rect 2411 6556 2475 6560
rect 2411 6500 2415 6556
rect 2415 6500 2471 6556
rect 2471 6500 2475 6556
rect 2411 6496 2475 6500
rect 2491 6556 2555 6560
rect 2491 6500 2495 6556
rect 2495 6500 2551 6556
rect 2551 6500 2555 6556
rect 2491 6496 2555 6500
rect 5953 6556 6017 6560
rect 5953 6500 5957 6556
rect 5957 6500 6013 6556
rect 6013 6500 6017 6556
rect 5953 6496 6017 6500
rect 6033 6556 6097 6560
rect 6033 6500 6037 6556
rect 6037 6500 6093 6556
rect 6093 6500 6097 6556
rect 6033 6496 6097 6500
rect 6113 6556 6177 6560
rect 6113 6500 6117 6556
rect 6117 6500 6173 6556
rect 6173 6500 6177 6556
rect 6113 6496 6177 6500
rect 6193 6556 6257 6560
rect 6193 6500 6197 6556
rect 6197 6500 6253 6556
rect 6253 6500 6257 6556
rect 6193 6496 6257 6500
rect 9655 6556 9719 6560
rect 9655 6500 9659 6556
rect 9659 6500 9715 6556
rect 9715 6500 9719 6556
rect 9655 6496 9719 6500
rect 9735 6556 9799 6560
rect 9735 6500 9739 6556
rect 9739 6500 9795 6556
rect 9795 6500 9799 6556
rect 9735 6496 9799 6500
rect 9815 6556 9879 6560
rect 9815 6500 9819 6556
rect 9819 6500 9875 6556
rect 9875 6500 9879 6556
rect 9815 6496 9879 6500
rect 9895 6556 9959 6560
rect 9895 6500 9899 6556
rect 9899 6500 9955 6556
rect 9955 6500 9959 6556
rect 9895 6496 9959 6500
rect 13357 6556 13421 6560
rect 13357 6500 13361 6556
rect 13361 6500 13417 6556
rect 13417 6500 13421 6556
rect 13357 6496 13421 6500
rect 13437 6556 13501 6560
rect 13437 6500 13441 6556
rect 13441 6500 13497 6556
rect 13497 6500 13501 6556
rect 13437 6496 13501 6500
rect 13517 6556 13581 6560
rect 13517 6500 13521 6556
rect 13521 6500 13577 6556
rect 13577 6500 13581 6556
rect 13517 6496 13581 6500
rect 13597 6556 13661 6560
rect 13597 6500 13601 6556
rect 13601 6500 13657 6556
rect 13657 6500 13661 6556
rect 13597 6496 13661 6500
rect 4102 6012 4166 6016
rect 4102 5956 4106 6012
rect 4106 5956 4162 6012
rect 4162 5956 4166 6012
rect 4102 5952 4166 5956
rect 4182 6012 4246 6016
rect 4182 5956 4186 6012
rect 4186 5956 4242 6012
rect 4242 5956 4246 6012
rect 4182 5952 4246 5956
rect 4262 6012 4326 6016
rect 4262 5956 4266 6012
rect 4266 5956 4322 6012
rect 4322 5956 4326 6012
rect 4262 5952 4326 5956
rect 4342 6012 4406 6016
rect 4342 5956 4346 6012
rect 4346 5956 4402 6012
rect 4402 5956 4406 6012
rect 4342 5952 4406 5956
rect 7804 6012 7868 6016
rect 7804 5956 7808 6012
rect 7808 5956 7864 6012
rect 7864 5956 7868 6012
rect 7804 5952 7868 5956
rect 7884 6012 7948 6016
rect 7884 5956 7888 6012
rect 7888 5956 7944 6012
rect 7944 5956 7948 6012
rect 7884 5952 7948 5956
rect 7964 6012 8028 6016
rect 7964 5956 7968 6012
rect 7968 5956 8024 6012
rect 8024 5956 8028 6012
rect 7964 5952 8028 5956
rect 8044 6012 8108 6016
rect 8044 5956 8048 6012
rect 8048 5956 8104 6012
rect 8104 5956 8108 6012
rect 8044 5952 8108 5956
rect 11506 6012 11570 6016
rect 11506 5956 11510 6012
rect 11510 5956 11566 6012
rect 11566 5956 11570 6012
rect 11506 5952 11570 5956
rect 11586 6012 11650 6016
rect 11586 5956 11590 6012
rect 11590 5956 11646 6012
rect 11646 5956 11650 6012
rect 11586 5952 11650 5956
rect 11666 6012 11730 6016
rect 11666 5956 11670 6012
rect 11670 5956 11726 6012
rect 11726 5956 11730 6012
rect 11666 5952 11730 5956
rect 11746 6012 11810 6016
rect 11746 5956 11750 6012
rect 11750 5956 11806 6012
rect 11806 5956 11810 6012
rect 11746 5952 11810 5956
rect 15208 6012 15272 6016
rect 15208 5956 15212 6012
rect 15212 5956 15268 6012
rect 15268 5956 15272 6012
rect 15208 5952 15272 5956
rect 15288 6012 15352 6016
rect 15288 5956 15292 6012
rect 15292 5956 15348 6012
rect 15348 5956 15352 6012
rect 15288 5952 15352 5956
rect 15368 6012 15432 6016
rect 15368 5956 15372 6012
rect 15372 5956 15428 6012
rect 15428 5956 15432 6012
rect 15368 5952 15432 5956
rect 15448 6012 15512 6016
rect 15448 5956 15452 6012
rect 15452 5956 15508 6012
rect 15508 5956 15512 6012
rect 15448 5952 15512 5956
rect 2251 5468 2315 5472
rect 2251 5412 2255 5468
rect 2255 5412 2311 5468
rect 2311 5412 2315 5468
rect 2251 5408 2315 5412
rect 2331 5468 2395 5472
rect 2331 5412 2335 5468
rect 2335 5412 2391 5468
rect 2391 5412 2395 5468
rect 2331 5408 2395 5412
rect 2411 5468 2475 5472
rect 2411 5412 2415 5468
rect 2415 5412 2471 5468
rect 2471 5412 2475 5468
rect 2411 5408 2475 5412
rect 2491 5468 2555 5472
rect 2491 5412 2495 5468
rect 2495 5412 2551 5468
rect 2551 5412 2555 5468
rect 2491 5408 2555 5412
rect 5953 5468 6017 5472
rect 5953 5412 5957 5468
rect 5957 5412 6013 5468
rect 6013 5412 6017 5468
rect 5953 5408 6017 5412
rect 6033 5468 6097 5472
rect 6033 5412 6037 5468
rect 6037 5412 6093 5468
rect 6093 5412 6097 5468
rect 6033 5408 6097 5412
rect 6113 5468 6177 5472
rect 6113 5412 6117 5468
rect 6117 5412 6173 5468
rect 6173 5412 6177 5468
rect 6113 5408 6177 5412
rect 6193 5468 6257 5472
rect 6193 5412 6197 5468
rect 6197 5412 6253 5468
rect 6253 5412 6257 5468
rect 6193 5408 6257 5412
rect 9655 5468 9719 5472
rect 9655 5412 9659 5468
rect 9659 5412 9715 5468
rect 9715 5412 9719 5468
rect 9655 5408 9719 5412
rect 9735 5468 9799 5472
rect 9735 5412 9739 5468
rect 9739 5412 9795 5468
rect 9795 5412 9799 5468
rect 9735 5408 9799 5412
rect 9815 5468 9879 5472
rect 9815 5412 9819 5468
rect 9819 5412 9875 5468
rect 9875 5412 9879 5468
rect 9815 5408 9879 5412
rect 9895 5468 9959 5472
rect 9895 5412 9899 5468
rect 9899 5412 9955 5468
rect 9955 5412 9959 5468
rect 9895 5408 9959 5412
rect 13357 5468 13421 5472
rect 13357 5412 13361 5468
rect 13361 5412 13417 5468
rect 13417 5412 13421 5468
rect 13357 5408 13421 5412
rect 13437 5468 13501 5472
rect 13437 5412 13441 5468
rect 13441 5412 13497 5468
rect 13497 5412 13501 5468
rect 13437 5408 13501 5412
rect 13517 5468 13581 5472
rect 13517 5412 13521 5468
rect 13521 5412 13577 5468
rect 13577 5412 13581 5468
rect 13517 5408 13581 5412
rect 13597 5468 13661 5472
rect 13597 5412 13601 5468
rect 13601 5412 13657 5468
rect 13657 5412 13661 5468
rect 13597 5408 13661 5412
rect 4102 4924 4166 4928
rect 4102 4868 4106 4924
rect 4106 4868 4162 4924
rect 4162 4868 4166 4924
rect 4102 4864 4166 4868
rect 4182 4924 4246 4928
rect 4182 4868 4186 4924
rect 4186 4868 4242 4924
rect 4242 4868 4246 4924
rect 4182 4864 4246 4868
rect 4262 4924 4326 4928
rect 4262 4868 4266 4924
rect 4266 4868 4322 4924
rect 4322 4868 4326 4924
rect 4262 4864 4326 4868
rect 4342 4924 4406 4928
rect 4342 4868 4346 4924
rect 4346 4868 4402 4924
rect 4402 4868 4406 4924
rect 4342 4864 4406 4868
rect 7804 4924 7868 4928
rect 7804 4868 7808 4924
rect 7808 4868 7864 4924
rect 7864 4868 7868 4924
rect 7804 4864 7868 4868
rect 7884 4924 7948 4928
rect 7884 4868 7888 4924
rect 7888 4868 7944 4924
rect 7944 4868 7948 4924
rect 7884 4864 7948 4868
rect 7964 4924 8028 4928
rect 7964 4868 7968 4924
rect 7968 4868 8024 4924
rect 8024 4868 8028 4924
rect 7964 4864 8028 4868
rect 8044 4924 8108 4928
rect 8044 4868 8048 4924
rect 8048 4868 8104 4924
rect 8104 4868 8108 4924
rect 8044 4864 8108 4868
rect 11506 4924 11570 4928
rect 11506 4868 11510 4924
rect 11510 4868 11566 4924
rect 11566 4868 11570 4924
rect 11506 4864 11570 4868
rect 11586 4924 11650 4928
rect 11586 4868 11590 4924
rect 11590 4868 11646 4924
rect 11646 4868 11650 4924
rect 11586 4864 11650 4868
rect 11666 4924 11730 4928
rect 11666 4868 11670 4924
rect 11670 4868 11726 4924
rect 11726 4868 11730 4924
rect 11666 4864 11730 4868
rect 11746 4924 11810 4928
rect 11746 4868 11750 4924
rect 11750 4868 11806 4924
rect 11806 4868 11810 4924
rect 11746 4864 11810 4868
rect 15208 4924 15272 4928
rect 15208 4868 15212 4924
rect 15212 4868 15268 4924
rect 15268 4868 15272 4924
rect 15208 4864 15272 4868
rect 15288 4924 15352 4928
rect 15288 4868 15292 4924
rect 15292 4868 15348 4924
rect 15348 4868 15352 4924
rect 15288 4864 15352 4868
rect 15368 4924 15432 4928
rect 15368 4868 15372 4924
rect 15372 4868 15428 4924
rect 15428 4868 15432 4924
rect 15368 4864 15432 4868
rect 15448 4924 15512 4928
rect 15448 4868 15452 4924
rect 15452 4868 15508 4924
rect 15508 4868 15512 4924
rect 15448 4864 15512 4868
rect 2251 4380 2315 4384
rect 2251 4324 2255 4380
rect 2255 4324 2311 4380
rect 2311 4324 2315 4380
rect 2251 4320 2315 4324
rect 2331 4380 2395 4384
rect 2331 4324 2335 4380
rect 2335 4324 2391 4380
rect 2391 4324 2395 4380
rect 2331 4320 2395 4324
rect 2411 4380 2475 4384
rect 2411 4324 2415 4380
rect 2415 4324 2471 4380
rect 2471 4324 2475 4380
rect 2411 4320 2475 4324
rect 2491 4380 2555 4384
rect 2491 4324 2495 4380
rect 2495 4324 2551 4380
rect 2551 4324 2555 4380
rect 2491 4320 2555 4324
rect 5953 4380 6017 4384
rect 5953 4324 5957 4380
rect 5957 4324 6013 4380
rect 6013 4324 6017 4380
rect 5953 4320 6017 4324
rect 6033 4380 6097 4384
rect 6033 4324 6037 4380
rect 6037 4324 6093 4380
rect 6093 4324 6097 4380
rect 6033 4320 6097 4324
rect 6113 4380 6177 4384
rect 6113 4324 6117 4380
rect 6117 4324 6173 4380
rect 6173 4324 6177 4380
rect 6113 4320 6177 4324
rect 6193 4380 6257 4384
rect 6193 4324 6197 4380
rect 6197 4324 6253 4380
rect 6253 4324 6257 4380
rect 6193 4320 6257 4324
rect 9655 4380 9719 4384
rect 9655 4324 9659 4380
rect 9659 4324 9715 4380
rect 9715 4324 9719 4380
rect 9655 4320 9719 4324
rect 9735 4380 9799 4384
rect 9735 4324 9739 4380
rect 9739 4324 9795 4380
rect 9795 4324 9799 4380
rect 9735 4320 9799 4324
rect 9815 4380 9879 4384
rect 9815 4324 9819 4380
rect 9819 4324 9875 4380
rect 9875 4324 9879 4380
rect 9815 4320 9879 4324
rect 9895 4380 9959 4384
rect 9895 4324 9899 4380
rect 9899 4324 9955 4380
rect 9955 4324 9959 4380
rect 9895 4320 9959 4324
rect 13357 4380 13421 4384
rect 13357 4324 13361 4380
rect 13361 4324 13417 4380
rect 13417 4324 13421 4380
rect 13357 4320 13421 4324
rect 13437 4380 13501 4384
rect 13437 4324 13441 4380
rect 13441 4324 13497 4380
rect 13497 4324 13501 4380
rect 13437 4320 13501 4324
rect 13517 4380 13581 4384
rect 13517 4324 13521 4380
rect 13521 4324 13577 4380
rect 13577 4324 13581 4380
rect 13517 4320 13581 4324
rect 13597 4380 13661 4384
rect 13597 4324 13601 4380
rect 13601 4324 13657 4380
rect 13657 4324 13661 4380
rect 13597 4320 13661 4324
rect 4102 3836 4166 3840
rect 4102 3780 4106 3836
rect 4106 3780 4162 3836
rect 4162 3780 4166 3836
rect 4102 3776 4166 3780
rect 4182 3836 4246 3840
rect 4182 3780 4186 3836
rect 4186 3780 4242 3836
rect 4242 3780 4246 3836
rect 4182 3776 4246 3780
rect 4262 3836 4326 3840
rect 4262 3780 4266 3836
rect 4266 3780 4322 3836
rect 4322 3780 4326 3836
rect 4262 3776 4326 3780
rect 4342 3836 4406 3840
rect 4342 3780 4346 3836
rect 4346 3780 4402 3836
rect 4402 3780 4406 3836
rect 4342 3776 4406 3780
rect 7804 3836 7868 3840
rect 7804 3780 7808 3836
rect 7808 3780 7864 3836
rect 7864 3780 7868 3836
rect 7804 3776 7868 3780
rect 7884 3836 7948 3840
rect 7884 3780 7888 3836
rect 7888 3780 7944 3836
rect 7944 3780 7948 3836
rect 7884 3776 7948 3780
rect 7964 3836 8028 3840
rect 7964 3780 7968 3836
rect 7968 3780 8024 3836
rect 8024 3780 8028 3836
rect 7964 3776 8028 3780
rect 8044 3836 8108 3840
rect 8044 3780 8048 3836
rect 8048 3780 8104 3836
rect 8104 3780 8108 3836
rect 8044 3776 8108 3780
rect 11506 3836 11570 3840
rect 11506 3780 11510 3836
rect 11510 3780 11566 3836
rect 11566 3780 11570 3836
rect 11506 3776 11570 3780
rect 11586 3836 11650 3840
rect 11586 3780 11590 3836
rect 11590 3780 11646 3836
rect 11646 3780 11650 3836
rect 11586 3776 11650 3780
rect 11666 3836 11730 3840
rect 11666 3780 11670 3836
rect 11670 3780 11726 3836
rect 11726 3780 11730 3836
rect 11666 3776 11730 3780
rect 11746 3836 11810 3840
rect 11746 3780 11750 3836
rect 11750 3780 11806 3836
rect 11806 3780 11810 3836
rect 11746 3776 11810 3780
rect 15208 3836 15272 3840
rect 15208 3780 15212 3836
rect 15212 3780 15268 3836
rect 15268 3780 15272 3836
rect 15208 3776 15272 3780
rect 15288 3836 15352 3840
rect 15288 3780 15292 3836
rect 15292 3780 15348 3836
rect 15348 3780 15352 3836
rect 15288 3776 15352 3780
rect 15368 3836 15432 3840
rect 15368 3780 15372 3836
rect 15372 3780 15428 3836
rect 15428 3780 15432 3836
rect 15368 3776 15432 3780
rect 15448 3836 15512 3840
rect 15448 3780 15452 3836
rect 15452 3780 15508 3836
rect 15508 3780 15512 3836
rect 15448 3776 15512 3780
rect 2251 3292 2315 3296
rect 2251 3236 2255 3292
rect 2255 3236 2311 3292
rect 2311 3236 2315 3292
rect 2251 3232 2315 3236
rect 2331 3292 2395 3296
rect 2331 3236 2335 3292
rect 2335 3236 2391 3292
rect 2391 3236 2395 3292
rect 2331 3232 2395 3236
rect 2411 3292 2475 3296
rect 2411 3236 2415 3292
rect 2415 3236 2471 3292
rect 2471 3236 2475 3292
rect 2411 3232 2475 3236
rect 2491 3292 2555 3296
rect 2491 3236 2495 3292
rect 2495 3236 2551 3292
rect 2551 3236 2555 3292
rect 2491 3232 2555 3236
rect 5953 3292 6017 3296
rect 5953 3236 5957 3292
rect 5957 3236 6013 3292
rect 6013 3236 6017 3292
rect 5953 3232 6017 3236
rect 6033 3292 6097 3296
rect 6033 3236 6037 3292
rect 6037 3236 6093 3292
rect 6093 3236 6097 3292
rect 6033 3232 6097 3236
rect 6113 3292 6177 3296
rect 6113 3236 6117 3292
rect 6117 3236 6173 3292
rect 6173 3236 6177 3292
rect 6113 3232 6177 3236
rect 6193 3292 6257 3296
rect 6193 3236 6197 3292
rect 6197 3236 6253 3292
rect 6253 3236 6257 3292
rect 6193 3232 6257 3236
rect 9655 3292 9719 3296
rect 9655 3236 9659 3292
rect 9659 3236 9715 3292
rect 9715 3236 9719 3292
rect 9655 3232 9719 3236
rect 9735 3292 9799 3296
rect 9735 3236 9739 3292
rect 9739 3236 9795 3292
rect 9795 3236 9799 3292
rect 9735 3232 9799 3236
rect 9815 3292 9879 3296
rect 9815 3236 9819 3292
rect 9819 3236 9875 3292
rect 9875 3236 9879 3292
rect 9815 3232 9879 3236
rect 9895 3292 9959 3296
rect 9895 3236 9899 3292
rect 9899 3236 9955 3292
rect 9955 3236 9959 3292
rect 9895 3232 9959 3236
rect 13357 3292 13421 3296
rect 13357 3236 13361 3292
rect 13361 3236 13417 3292
rect 13417 3236 13421 3292
rect 13357 3232 13421 3236
rect 13437 3292 13501 3296
rect 13437 3236 13441 3292
rect 13441 3236 13497 3292
rect 13497 3236 13501 3292
rect 13437 3232 13501 3236
rect 13517 3292 13581 3296
rect 13517 3236 13521 3292
rect 13521 3236 13577 3292
rect 13577 3236 13581 3292
rect 13517 3232 13581 3236
rect 13597 3292 13661 3296
rect 13597 3236 13601 3292
rect 13601 3236 13657 3292
rect 13657 3236 13661 3292
rect 13597 3232 13661 3236
rect 4102 2748 4166 2752
rect 4102 2692 4106 2748
rect 4106 2692 4162 2748
rect 4162 2692 4166 2748
rect 4102 2688 4166 2692
rect 4182 2748 4246 2752
rect 4182 2692 4186 2748
rect 4186 2692 4242 2748
rect 4242 2692 4246 2748
rect 4182 2688 4246 2692
rect 4262 2748 4326 2752
rect 4262 2692 4266 2748
rect 4266 2692 4322 2748
rect 4322 2692 4326 2748
rect 4262 2688 4326 2692
rect 4342 2748 4406 2752
rect 4342 2692 4346 2748
rect 4346 2692 4402 2748
rect 4402 2692 4406 2748
rect 4342 2688 4406 2692
rect 7804 2748 7868 2752
rect 7804 2692 7808 2748
rect 7808 2692 7864 2748
rect 7864 2692 7868 2748
rect 7804 2688 7868 2692
rect 7884 2748 7948 2752
rect 7884 2692 7888 2748
rect 7888 2692 7944 2748
rect 7944 2692 7948 2748
rect 7884 2688 7948 2692
rect 7964 2748 8028 2752
rect 7964 2692 7968 2748
rect 7968 2692 8024 2748
rect 8024 2692 8028 2748
rect 7964 2688 8028 2692
rect 8044 2748 8108 2752
rect 8044 2692 8048 2748
rect 8048 2692 8104 2748
rect 8104 2692 8108 2748
rect 8044 2688 8108 2692
rect 11506 2748 11570 2752
rect 11506 2692 11510 2748
rect 11510 2692 11566 2748
rect 11566 2692 11570 2748
rect 11506 2688 11570 2692
rect 11586 2748 11650 2752
rect 11586 2692 11590 2748
rect 11590 2692 11646 2748
rect 11646 2692 11650 2748
rect 11586 2688 11650 2692
rect 11666 2748 11730 2752
rect 11666 2692 11670 2748
rect 11670 2692 11726 2748
rect 11726 2692 11730 2748
rect 11666 2688 11730 2692
rect 11746 2748 11810 2752
rect 11746 2692 11750 2748
rect 11750 2692 11806 2748
rect 11806 2692 11810 2748
rect 11746 2688 11810 2692
rect 15208 2748 15272 2752
rect 15208 2692 15212 2748
rect 15212 2692 15268 2748
rect 15268 2692 15272 2748
rect 15208 2688 15272 2692
rect 15288 2748 15352 2752
rect 15288 2692 15292 2748
rect 15292 2692 15348 2748
rect 15348 2692 15352 2748
rect 15288 2688 15352 2692
rect 15368 2748 15432 2752
rect 15368 2692 15372 2748
rect 15372 2692 15428 2748
rect 15428 2692 15432 2748
rect 15368 2688 15432 2692
rect 15448 2748 15512 2752
rect 15448 2692 15452 2748
rect 15452 2692 15508 2748
rect 15508 2692 15512 2748
rect 15448 2688 15512 2692
rect 2251 2204 2315 2208
rect 2251 2148 2255 2204
rect 2255 2148 2311 2204
rect 2311 2148 2315 2204
rect 2251 2144 2315 2148
rect 2331 2204 2395 2208
rect 2331 2148 2335 2204
rect 2335 2148 2391 2204
rect 2391 2148 2395 2204
rect 2331 2144 2395 2148
rect 2411 2204 2475 2208
rect 2411 2148 2415 2204
rect 2415 2148 2471 2204
rect 2471 2148 2475 2204
rect 2411 2144 2475 2148
rect 2491 2204 2555 2208
rect 2491 2148 2495 2204
rect 2495 2148 2551 2204
rect 2551 2148 2555 2204
rect 2491 2144 2555 2148
rect 5953 2204 6017 2208
rect 5953 2148 5957 2204
rect 5957 2148 6013 2204
rect 6013 2148 6017 2204
rect 5953 2144 6017 2148
rect 6033 2204 6097 2208
rect 6033 2148 6037 2204
rect 6037 2148 6093 2204
rect 6093 2148 6097 2204
rect 6033 2144 6097 2148
rect 6113 2204 6177 2208
rect 6113 2148 6117 2204
rect 6117 2148 6173 2204
rect 6173 2148 6177 2204
rect 6113 2144 6177 2148
rect 6193 2204 6257 2208
rect 6193 2148 6197 2204
rect 6197 2148 6253 2204
rect 6253 2148 6257 2204
rect 6193 2144 6257 2148
rect 9655 2204 9719 2208
rect 9655 2148 9659 2204
rect 9659 2148 9715 2204
rect 9715 2148 9719 2204
rect 9655 2144 9719 2148
rect 9735 2204 9799 2208
rect 9735 2148 9739 2204
rect 9739 2148 9795 2204
rect 9795 2148 9799 2204
rect 9735 2144 9799 2148
rect 9815 2204 9879 2208
rect 9815 2148 9819 2204
rect 9819 2148 9875 2204
rect 9875 2148 9879 2204
rect 9815 2144 9879 2148
rect 9895 2204 9959 2208
rect 9895 2148 9899 2204
rect 9899 2148 9955 2204
rect 9955 2148 9959 2204
rect 9895 2144 9959 2148
rect 13357 2204 13421 2208
rect 13357 2148 13361 2204
rect 13361 2148 13417 2204
rect 13417 2148 13421 2204
rect 13357 2144 13421 2148
rect 13437 2204 13501 2208
rect 13437 2148 13441 2204
rect 13441 2148 13497 2204
rect 13497 2148 13501 2204
rect 13437 2144 13501 2148
rect 13517 2204 13581 2208
rect 13517 2148 13521 2204
rect 13521 2148 13577 2204
rect 13577 2148 13581 2204
rect 13517 2144 13581 2148
rect 13597 2204 13661 2208
rect 13597 2148 13601 2204
rect 13601 2148 13657 2204
rect 13657 2148 13661 2204
rect 13597 2144 13661 2148
rect 4102 1660 4166 1664
rect 4102 1604 4106 1660
rect 4106 1604 4162 1660
rect 4162 1604 4166 1660
rect 4102 1600 4166 1604
rect 4182 1660 4246 1664
rect 4182 1604 4186 1660
rect 4186 1604 4242 1660
rect 4242 1604 4246 1660
rect 4182 1600 4246 1604
rect 4262 1660 4326 1664
rect 4262 1604 4266 1660
rect 4266 1604 4322 1660
rect 4322 1604 4326 1660
rect 4262 1600 4326 1604
rect 4342 1660 4406 1664
rect 4342 1604 4346 1660
rect 4346 1604 4402 1660
rect 4402 1604 4406 1660
rect 4342 1600 4406 1604
rect 7804 1660 7868 1664
rect 7804 1604 7808 1660
rect 7808 1604 7864 1660
rect 7864 1604 7868 1660
rect 7804 1600 7868 1604
rect 7884 1660 7948 1664
rect 7884 1604 7888 1660
rect 7888 1604 7944 1660
rect 7944 1604 7948 1660
rect 7884 1600 7948 1604
rect 7964 1660 8028 1664
rect 7964 1604 7968 1660
rect 7968 1604 8024 1660
rect 8024 1604 8028 1660
rect 7964 1600 8028 1604
rect 8044 1660 8108 1664
rect 8044 1604 8048 1660
rect 8048 1604 8104 1660
rect 8104 1604 8108 1660
rect 8044 1600 8108 1604
rect 11506 1660 11570 1664
rect 11506 1604 11510 1660
rect 11510 1604 11566 1660
rect 11566 1604 11570 1660
rect 11506 1600 11570 1604
rect 11586 1660 11650 1664
rect 11586 1604 11590 1660
rect 11590 1604 11646 1660
rect 11646 1604 11650 1660
rect 11586 1600 11650 1604
rect 11666 1660 11730 1664
rect 11666 1604 11670 1660
rect 11670 1604 11726 1660
rect 11726 1604 11730 1660
rect 11666 1600 11730 1604
rect 11746 1660 11810 1664
rect 11746 1604 11750 1660
rect 11750 1604 11806 1660
rect 11806 1604 11810 1660
rect 11746 1600 11810 1604
rect 15208 1660 15272 1664
rect 15208 1604 15212 1660
rect 15212 1604 15268 1660
rect 15268 1604 15272 1660
rect 15208 1600 15272 1604
rect 15288 1660 15352 1664
rect 15288 1604 15292 1660
rect 15292 1604 15348 1660
rect 15348 1604 15352 1660
rect 15288 1600 15352 1604
rect 15368 1660 15432 1664
rect 15368 1604 15372 1660
rect 15372 1604 15428 1660
rect 15428 1604 15432 1660
rect 15368 1600 15432 1604
rect 15448 1660 15512 1664
rect 15448 1604 15452 1660
rect 15452 1604 15508 1660
rect 15508 1604 15512 1660
rect 15448 1600 15512 1604
rect 2251 1116 2315 1120
rect 2251 1060 2255 1116
rect 2255 1060 2311 1116
rect 2311 1060 2315 1116
rect 2251 1056 2315 1060
rect 2331 1116 2395 1120
rect 2331 1060 2335 1116
rect 2335 1060 2391 1116
rect 2391 1060 2395 1116
rect 2331 1056 2395 1060
rect 2411 1116 2475 1120
rect 2411 1060 2415 1116
rect 2415 1060 2471 1116
rect 2471 1060 2475 1116
rect 2411 1056 2475 1060
rect 2491 1116 2555 1120
rect 2491 1060 2495 1116
rect 2495 1060 2551 1116
rect 2551 1060 2555 1116
rect 2491 1056 2555 1060
rect 5953 1116 6017 1120
rect 5953 1060 5957 1116
rect 5957 1060 6013 1116
rect 6013 1060 6017 1116
rect 5953 1056 6017 1060
rect 6033 1116 6097 1120
rect 6033 1060 6037 1116
rect 6037 1060 6093 1116
rect 6093 1060 6097 1116
rect 6033 1056 6097 1060
rect 6113 1116 6177 1120
rect 6113 1060 6117 1116
rect 6117 1060 6173 1116
rect 6173 1060 6177 1116
rect 6113 1056 6177 1060
rect 6193 1116 6257 1120
rect 6193 1060 6197 1116
rect 6197 1060 6253 1116
rect 6253 1060 6257 1116
rect 6193 1056 6257 1060
rect 9655 1116 9719 1120
rect 9655 1060 9659 1116
rect 9659 1060 9715 1116
rect 9715 1060 9719 1116
rect 9655 1056 9719 1060
rect 9735 1116 9799 1120
rect 9735 1060 9739 1116
rect 9739 1060 9795 1116
rect 9795 1060 9799 1116
rect 9735 1056 9799 1060
rect 9815 1116 9879 1120
rect 9815 1060 9819 1116
rect 9819 1060 9875 1116
rect 9875 1060 9879 1116
rect 9815 1056 9879 1060
rect 9895 1116 9959 1120
rect 9895 1060 9899 1116
rect 9899 1060 9955 1116
rect 9955 1060 9959 1116
rect 9895 1056 9959 1060
rect 13357 1116 13421 1120
rect 13357 1060 13361 1116
rect 13361 1060 13417 1116
rect 13417 1060 13421 1116
rect 13357 1056 13421 1060
rect 13437 1116 13501 1120
rect 13437 1060 13441 1116
rect 13441 1060 13497 1116
rect 13497 1060 13501 1116
rect 13437 1056 13501 1060
rect 13517 1116 13581 1120
rect 13517 1060 13521 1116
rect 13521 1060 13577 1116
rect 13577 1060 13581 1116
rect 13517 1056 13581 1060
rect 13597 1116 13661 1120
rect 13597 1060 13601 1116
rect 13601 1060 13657 1116
rect 13657 1060 13661 1116
rect 13597 1056 13661 1060
rect 4102 572 4166 576
rect 4102 516 4106 572
rect 4106 516 4162 572
rect 4162 516 4166 572
rect 4102 512 4166 516
rect 4182 572 4246 576
rect 4182 516 4186 572
rect 4186 516 4242 572
rect 4242 516 4246 572
rect 4182 512 4246 516
rect 4262 572 4326 576
rect 4262 516 4266 572
rect 4266 516 4322 572
rect 4322 516 4326 572
rect 4262 512 4326 516
rect 4342 572 4406 576
rect 4342 516 4346 572
rect 4346 516 4402 572
rect 4402 516 4406 572
rect 4342 512 4406 516
rect 7804 572 7868 576
rect 7804 516 7808 572
rect 7808 516 7864 572
rect 7864 516 7868 572
rect 7804 512 7868 516
rect 7884 572 7948 576
rect 7884 516 7888 572
rect 7888 516 7944 572
rect 7944 516 7948 572
rect 7884 512 7948 516
rect 7964 572 8028 576
rect 7964 516 7968 572
rect 7968 516 8024 572
rect 8024 516 8028 572
rect 7964 512 8028 516
rect 8044 572 8108 576
rect 8044 516 8048 572
rect 8048 516 8104 572
rect 8104 516 8108 572
rect 8044 512 8108 516
rect 11506 572 11570 576
rect 11506 516 11510 572
rect 11510 516 11566 572
rect 11566 516 11570 572
rect 11506 512 11570 516
rect 11586 572 11650 576
rect 11586 516 11590 572
rect 11590 516 11646 572
rect 11646 516 11650 572
rect 11586 512 11650 516
rect 11666 572 11730 576
rect 11666 516 11670 572
rect 11670 516 11726 572
rect 11726 516 11730 572
rect 11666 512 11730 516
rect 11746 572 11810 576
rect 11746 516 11750 572
rect 11750 516 11806 572
rect 11806 516 11810 572
rect 11746 512 11810 516
rect 15208 572 15272 576
rect 15208 516 15212 572
rect 15212 516 15268 572
rect 15268 516 15272 572
rect 15208 512 15272 516
rect 15288 572 15352 576
rect 15288 516 15292 572
rect 15292 516 15348 572
rect 15348 516 15352 572
rect 15288 512 15352 516
rect 15368 572 15432 576
rect 15368 516 15372 572
rect 15372 516 15428 572
rect 15428 516 15432 572
rect 15368 512 15432 516
rect 15448 572 15512 576
rect 15448 516 15452 572
rect 15452 516 15508 572
rect 15508 516 15512 572
rect 15448 512 15512 516
<< metal4 >>
rect 2243 15264 2563 15280
rect 2243 15200 2251 15264
rect 2315 15200 2331 15264
rect 2395 15200 2411 15264
rect 2475 15200 2491 15264
rect 2555 15200 2563 15264
rect 2243 14176 2563 15200
rect 2243 14112 2251 14176
rect 2315 14112 2331 14176
rect 2395 14112 2411 14176
rect 2475 14112 2491 14176
rect 2555 14112 2563 14176
rect 2243 13088 2563 14112
rect 2243 13024 2251 13088
rect 2315 13024 2331 13088
rect 2395 13024 2411 13088
rect 2475 13024 2491 13088
rect 2555 13024 2563 13088
rect 2243 12000 2563 13024
rect 2243 11936 2251 12000
rect 2315 11936 2331 12000
rect 2395 11936 2411 12000
rect 2475 11936 2491 12000
rect 2555 11936 2563 12000
rect 2243 10912 2563 11936
rect 2243 10848 2251 10912
rect 2315 10848 2331 10912
rect 2395 10848 2411 10912
rect 2475 10848 2491 10912
rect 2555 10848 2563 10912
rect 2243 9824 2563 10848
rect 2243 9760 2251 9824
rect 2315 9760 2331 9824
rect 2395 9760 2411 9824
rect 2475 9760 2491 9824
rect 2555 9760 2563 9824
rect 2243 8736 2563 9760
rect 2243 8672 2251 8736
rect 2315 8672 2331 8736
rect 2395 8672 2411 8736
rect 2475 8672 2491 8736
rect 2555 8672 2563 8736
rect 2243 7648 2563 8672
rect 2243 7584 2251 7648
rect 2315 7584 2331 7648
rect 2395 7584 2411 7648
rect 2475 7584 2491 7648
rect 2555 7584 2563 7648
rect 2243 6560 2563 7584
rect 2243 6496 2251 6560
rect 2315 6496 2331 6560
rect 2395 6496 2411 6560
rect 2475 6496 2491 6560
rect 2555 6496 2563 6560
rect 2243 5472 2563 6496
rect 2243 5408 2251 5472
rect 2315 5408 2331 5472
rect 2395 5408 2411 5472
rect 2475 5408 2491 5472
rect 2555 5408 2563 5472
rect 2243 4384 2563 5408
rect 2243 4320 2251 4384
rect 2315 4320 2331 4384
rect 2395 4320 2411 4384
rect 2475 4320 2491 4384
rect 2555 4320 2563 4384
rect 2243 3296 2563 4320
rect 2243 3232 2251 3296
rect 2315 3232 2331 3296
rect 2395 3232 2411 3296
rect 2475 3232 2491 3296
rect 2555 3232 2563 3296
rect 2243 2208 2563 3232
rect 2243 2144 2251 2208
rect 2315 2144 2331 2208
rect 2395 2144 2411 2208
rect 2475 2144 2491 2208
rect 2555 2144 2563 2208
rect 2243 1120 2563 2144
rect 2243 1056 2251 1120
rect 2315 1056 2331 1120
rect 2395 1056 2411 1120
rect 2475 1056 2491 1120
rect 2555 1056 2563 1120
rect 2243 496 2563 1056
rect 4094 14720 4414 15280
rect 4094 14656 4102 14720
rect 4166 14656 4182 14720
rect 4246 14656 4262 14720
rect 4326 14656 4342 14720
rect 4406 14656 4414 14720
rect 4094 13632 4414 14656
rect 4094 13568 4102 13632
rect 4166 13568 4182 13632
rect 4246 13568 4262 13632
rect 4326 13568 4342 13632
rect 4406 13568 4414 13632
rect 4094 12544 4414 13568
rect 4094 12480 4102 12544
rect 4166 12480 4182 12544
rect 4246 12480 4262 12544
rect 4326 12480 4342 12544
rect 4406 12480 4414 12544
rect 4094 11456 4414 12480
rect 4094 11392 4102 11456
rect 4166 11392 4182 11456
rect 4246 11392 4262 11456
rect 4326 11392 4342 11456
rect 4406 11392 4414 11456
rect 4094 10368 4414 11392
rect 4094 10304 4102 10368
rect 4166 10304 4182 10368
rect 4246 10304 4262 10368
rect 4326 10304 4342 10368
rect 4406 10304 4414 10368
rect 4094 9280 4414 10304
rect 4094 9216 4102 9280
rect 4166 9216 4182 9280
rect 4246 9216 4262 9280
rect 4326 9216 4342 9280
rect 4406 9216 4414 9280
rect 4094 8192 4414 9216
rect 4094 8128 4102 8192
rect 4166 8128 4182 8192
rect 4246 8128 4262 8192
rect 4326 8128 4342 8192
rect 4406 8128 4414 8192
rect 4094 7104 4414 8128
rect 4094 7040 4102 7104
rect 4166 7040 4182 7104
rect 4246 7040 4262 7104
rect 4326 7040 4342 7104
rect 4406 7040 4414 7104
rect 4094 6016 4414 7040
rect 4094 5952 4102 6016
rect 4166 5952 4182 6016
rect 4246 5952 4262 6016
rect 4326 5952 4342 6016
rect 4406 5952 4414 6016
rect 4094 4928 4414 5952
rect 4094 4864 4102 4928
rect 4166 4864 4182 4928
rect 4246 4864 4262 4928
rect 4326 4864 4342 4928
rect 4406 4864 4414 4928
rect 4094 3840 4414 4864
rect 4094 3776 4102 3840
rect 4166 3776 4182 3840
rect 4246 3776 4262 3840
rect 4326 3776 4342 3840
rect 4406 3776 4414 3840
rect 4094 2752 4414 3776
rect 4094 2688 4102 2752
rect 4166 2688 4182 2752
rect 4246 2688 4262 2752
rect 4326 2688 4342 2752
rect 4406 2688 4414 2752
rect 4094 1664 4414 2688
rect 4094 1600 4102 1664
rect 4166 1600 4182 1664
rect 4246 1600 4262 1664
rect 4326 1600 4342 1664
rect 4406 1600 4414 1664
rect 4094 576 4414 1600
rect 4094 512 4102 576
rect 4166 512 4182 576
rect 4246 512 4262 576
rect 4326 512 4342 576
rect 4406 512 4414 576
rect 4094 496 4414 512
rect 5945 15264 6265 15280
rect 5945 15200 5953 15264
rect 6017 15200 6033 15264
rect 6097 15200 6113 15264
rect 6177 15200 6193 15264
rect 6257 15200 6265 15264
rect 5945 14176 6265 15200
rect 5945 14112 5953 14176
rect 6017 14112 6033 14176
rect 6097 14112 6113 14176
rect 6177 14112 6193 14176
rect 6257 14112 6265 14176
rect 5945 13088 6265 14112
rect 5945 13024 5953 13088
rect 6017 13024 6033 13088
rect 6097 13024 6113 13088
rect 6177 13024 6193 13088
rect 6257 13024 6265 13088
rect 5945 12000 6265 13024
rect 5945 11936 5953 12000
rect 6017 11936 6033 12000
rect 6097 11936 6113 12000
rect 6177 11936 6193 12000
rect 6257 11936 6265 12000
rect 5945 10912 6265 11936
rect 5945 10848 5953 10912
rect 6017 10848 6033 10912
rect 6097 10848 6113 10912
rect 6177 10848 6193 10912
rect 6257 10848 6265 10912
rect 5945 9824 6265 10848
rect 5945 9760 5953 9824
rect 6017 9760 6033 9824
rect 6097 9760 6113 9824
rect 6177 9760 6193 9824
rect 6257 9760 6265 9824
rect 5945 8736 6265 9760
rect 5945 8672 5953 8736
rect 6017 8672 6033 8736
rect 6097 8672 6113 8736
rect 6177 8672 6193 8736
rect 6257 8672 6265 8736
rect 5945 7648 6265 8672
rect 5945 7584 5953 7648
rect 6017 7584 6033 7648
rect 6097 7584 6113 7648
rect 6177 7584 6193 7648
rect 6257 7584 6265 7648
rect 5945 6560 6265 7584
rect 5945 6496 5953 6560
rect 6017 6496 6033 6560
rect 6097 6496 6113 6560
rect 6177 6496 6193 6560
rect 6257 6496 6265 6560
rect 5945 5472 6265 6496
rect 5945 5408 5953 5472
rect 6017 5408 6033 5472
rect 6097 5408 6113 5472
rect 6177 5408 6193 5472
rect 6257 5408 6265 5472
rect 5945 4384 6265 5408
rect 5945 4320 5953 4384
rect 6017 4320 6033 4384
rect 6097 4320 6113 4384
rect 6177 4320 6193 4384
rect 6257 4320 6265 4384
rect 5945 3296 6265 4320
rect 5945 3232 5953 3296
rect 6017 3232 6033 3296
rect 6097 3232 6113 3296
rect 6177 3232 6193 3296
rect 6257 3232 6265 3296
rect 5945 2208 6265 3232
rect 5945 2144 5953 2208
rect 6017 2144 6033 2208
rect 6097 2144 6113 2208
rect 6177 2144 6193 2208
rect 6257 2144 6265 2208
rect 5945 1120 6265 2144
rect 5945 1056 5953 1120
rect 6017 1056 6033 1120
rect 6097 1056 6113 1120
rect 6177 1056 6193 1120
rect 6257 1056 6265 1120
rect 5945 496 6265 1056
rect 7796 14720 8116 15280
rect 7796 14656 7804 14720
rect 7868 14656 7884 14720
rect 7948 14656 7964 14720
rect 8028 14656 8044 14720
rect 8108 14656 8116 14720
rect 7796 13632 8116 14656
rect 7796 13568 7804 13632
rect 7868 13568 7884 13632
rect 7948 13568 7964 13632
rect 8028 13568 8044 13632
rect 8108 13568 8116 13632
rect 7796 12544 8116 13568
rect 7796 12480 7804 12544
rect 7868 12480 7884 12544
rect 7948 12480 7964 12544
rect 8028 12480 8044 12544
rect 8108 12480 8116 12544
rect 7796 11456 8116 12480
rect 7796 11392 7804 11456
rect 7868 11392 7884 11456
rect 7948 11392 7964 11456
rect 8028 11392 8044 11456
rect 8108 11392 8116 11456
rect 7796 10368 8116 11392
rect 7796 10304 7804 10368
rect 7868 10304 7884 10368
rect 7948 10304 7964 10368
rect 8028 10304 8044 10368
rect 8108 10304 8116 10368
rect 7796 9280 8116 10304
rect 7796 9216 7804 9280
rect 7868 9216 7884 9280
rect 7948 9216 7964 9280
rect 8028 9216 8044 9280
rect 8108 9216 8116 9280
rect 7796 8192 8116 9216
rect 7796 8128 7804 8192
rect 7868 8128 7884 8192
rect 7948 8128 7964 8192
rect 8028 8128 8044 8192
rect 8108 8128 8116 8192
rect 7796 7104 8116 8128
rect 7796 7040 7804 7104
rect 7868 7040 7884 7104
rect 7948 7040 7964 7104
rect 8028 7040 8044 7104
rect 8108 7040 8116 7104
rect 7796 6016 8116 7040
rect 7796 5952 7804 6016
rect 7868 5952 7884 6016
rect 7948 5952 7964 6016
rect 8028 5952 8044 6016
rect 8108 5952 8116 6016
rect 7796 4928 8116 5952
rect 7796 4864 7804 4928
rect 7868 4864 7884 4928
rect 7948 4864 7964 4928
rect 8028 4864 8044 4928
rect 8108 4864 8116 4928
rect 7796 3840 8116 4864
rect 7796 3776 7804 3840
rect 7868 3776 7884 3840
rect 7948 3776 7964 3840
rect 8028 3776 8044 3840
rect 8108 3776 8116 3840
rect 7796 2752 8116 3776
rect 7796 2688 7804 2752
rect 7868 2688 7884 2752
rect 7948 2688 7964 2752
rect 8028 2688 8044 2752
rect 8108 2688 8116 2752
rect 7796 1664 8116 2688
rect 7796 1600 7804 1664
rect 7868 1600 7884 1664
rect 7948 1600 7964 1664
rect 8028 1600 8044 1664
rect 8108 1600 8116 1664
rect 7796 576 8116 1600
rect 7796 512 7804 576
rect 7868 512 7884 576
rect 7948 512 7964 576
rect 8028 512 8044 576
rect 8108 512 8116 576
rect 7796 496 8116 512
rect 9647 15264 9967 15280
rect 9647 15200 9655 15264
rect 9719 15200 9735 15264
rect 9799 15200 9815 15264
rect 9879 15200 9895 15264
rect 9959 15200 9967 15264
rect 9647 14176 9967 15200
rect 9647 14112 9655 14176
rect 9719 14112 9735 14176
rect 9799 14112 9815 14176
rect 9879 14112 9895 14176
rect 9959 14112 9967 14176
rect 9647 13088 9967 14112
rect 9647 13024 9655 13088
rect 9719 13024 9735 13088
rect 9799 13024 9815 13088
rect 9879 13024 9895 13088
rect 9959 13024 9967 13088
rect 9647 12000 9967 13024
rect 9647 11936 9655 12000
rect 9719 11936 9735 12000
rect 9799 11936 9815 12000
rect 9879 11936 9895 12000
rect 9959 11936 9967 12000
rect 9647 10912 9967 11936
rect 9647 10848 9655 10912
rect 9719 10848 9735 10912
rect 9799 10848 9815 10912
rect 9879 10848 9895 10912
rect 9959 10848 9967 10912
rect 9647 9824 9967 10848
rect 9647 9760 9655 9824
rect 9719 9760 9735 9824
rect 9799 9760 9815 9824
rect 9879 9760 9895 9824
rect 9959 9760 9967 9824
rect 9647 8736 9967 9760
rect 9647 8672 9655 8736
rect 9719 8672 9735 8736
rect 9799 8672 9815 8736
rect 9879 8672 9895 8736
rect 9959 8672 9967 8736
rect 9647 7648 9967 8672
rect 9647 7584 9655 7648
rect 9719 7584 9735 7648
rect 9799 7584 9815 7648
rect 9879 7584 9895 7648
rect 9959 7584 9967 7648
rect 9647 6560 9967 7584
rect 9647 6496 9655 6560
rect 9719 6496 9735 6560
rect 9799 6496 9815 6560
rect 9879 6496 9895 6560
rect 9959 6496 9967 6560
rect 9647 5472 9967 6496
rect 9647 5408 9655 5472
rect 9719 5408 9735 5472
rect 9799 5408 9815 5472
rect 9879 5408 9895 5472
rect 9959 5408 9967 5472
rect 9647 4384 9967 5408
rect 9647 4320 9655 4384
rect 9719 4320 9735 4384
rect 9799 4320 9815 4384
rect 9879 4320 9895 4384
rect 9959 4320 9967 4384
rect 9647 3296 9967 4320
rect 9647 3232 9655 3296
rect 9719 3232 9735 3296
rect 9799 3232 9815 3296
rect 9879 3232 9895 3296
rect 9959 3232 9967 3296
rect 9647 2208 9967 3232
rect 9647 2144 9655 2208
rect 9719 2144 9735 2208
rect 9799 2144 9815 2208
rect 9879 2144 9895 2208
rect 9959 2144 9967 2208
rect 9647 1120 9967 2144
rect 9647 1056 9655 1120
rect 9719 1056 9735 1120
rect 9799 1056 9815 1120
rect 9879 1056 9895 1120
rect 9959 1056 9967 1120
rect 9647 496 9967 1056
rect 11498 14720 11818 15280
rect 11498 14656 11506 14720
rect 11570 14656 11586 14720
rect 11650 14656 11666 14720
rect 11730 14656 11746 14720
rect 11810 14656 11818 14720
rect 11498 13632 11818 14656
rect 11498 13568 11506 13632
rect 11570 13568 11586 13632
rect 11650 13568 11666 13632
rect 11730 13568 11746 13632
rect 11810 13568 11818 13632
rect 11498 12544 11818 13568
rect 11498 12480 11506 12544
rect 11570 12480 11586 12544
rect 11650 12480 11666 12544
rect 11730 12480 11746 12544
rect 11810 12480 11818 12544
rect 11498 11456 11818 12480
rect 11498 11392 11506 11456
rect 11570 11392 11586 11456
rect 11650 11392 11666 11456
rect 11730 11392 11746 11456
rect 11810 11392 11818 11456
rect 11498 10368 11818 11392
rect 11498 10304 11506 10368
rect 11570 10304 11586 10368
rect 11650 10304 11666 10368
rect 11730 10304 11746 10368
rect 11810 10304 11818 10368
rect 11498 9280 11818 10304
rect 11498 9216 11506 9280
rect 11570 9216 11586 9280
rect 11650 9216 11666 9280
rect 11730 9216 11746 9280
rect 11810 9216 11818 9280
rect 11498 8192 11818 9216
rect 11498 8128 11506 8192
rect 11570 8128 11586 8192
rect 11650 8128 11666 8192
rect 11730 8128 11746 8192
rect 11810 8128 11818 8192
rect 11498 7104 11818 8128
rect 11498 7040 11506 7104
rect 11570 7040 11586 7104
rect 11650 7040 11666 7104
rect 11730 7040 11746 7104
rect 11810 7040 11818 7104
rect 11498 6016 11818 7040
rect 11498 5952 11506 6016
rect 11570 5952 11586 6016
rect 11650 5952 11666 6016
rect 11730 5952 11746 6016
rect 11810 5952 11818 6016
rect 11498 4928 11818 5952
rect 11498 4864 11506 4928
rect 11570 4864 11586 4928
rect 11650 4864 11666 4928
rect 11730 4864 11746 4928
rect 11810 4864 11818 4928
rect 11498 3840 11818 4864
rect 11498 3776 11506 3840
rect 11570 3776 11586 3840
rect 11650 3776 11666 3840
rect 11730 3776 11746 3840
rect 11810 3776 11818 3840
rect 11498 2752 11818 3776
rect 11498 2688 11506 2752
rect 11570 2688 11586 2752
rect 11650 2688 11666 2752
rect 11730 2688 11746 2752
rect 11810 2688 11818 2752
rect 11498 1664 11818 2688
rect 11498 1600 11506 1664
rect 11570 1600 11586 1664
rect 11650 1600 11666 1664
rect 11730 1600 11746 1664
rect 11810 1600 11818 1664
rect 11498 576 11818 1600
rect 11498 512 11506 576
rect 11570 512 11586 576
rect 11650 512 11666 576
rect 11730 512 11746 576
rect 11810 512 11818 576
rect 11498 496 11818 512
rect 13349 15264 13669 15280
rect 13349 15200 13357 15264
rect 13421 15200 13437 15264
rect 13501 15200 13517 15264
rect 13581 15200 13597 15264
rect 13661 15200 13669 15264
rect 13349 14176 13669 15200
rect 13349 14112 13357 14176
rect 13421 14112 13437 14176
rect 13501 14112 13517 14176
rect 13581 14112 13597 14176
rect 13661 14112 13669 14176
rect 13349 13088 13669 14112
rect 13349 13024 13357 13088
rect 13421 13024 13437 13088
rect 13501 13024 13517 13088
rect 13581 13024 13597 13088
rect 13661 13024 13669 13088
rect 13349 12000 13669 13024
rect 13349 11936 13357 12000
rect 13421 11936 13437 12000
rect 13501 11936 13517 12000
rect 13581 11936 13597 12000
rect 13661 11936 13669 12000
rect 13349 10912 13669 11936
rect 13349 10848 13357 10912
rect 13421 10848 13437 10912
rect 13501 10848 13517 10912
rect 13581 10848 13597 10912
rect 13661 10848 13669 10912
rect 13349 9824 13669 10848
rect 13349 9760 13357 9824
rect 13421 9760 13437 9824
rect 13501 9760 13517 9824
rect 13581 9760 13597 9824
rect 13661 9760 13669 9824
rect 13349 8736 13669 9760
rect 13349 8672 13357 8736
rect 13421 8672 13437 8736
rect 13501 8672 13517 8736
rect 13581 8672 13597 8736
rect 13661 8672 13669 8736
rect 13349 7648 13669 8672
rect 13349 7584 13357 7648
rect 13421 7584 13437 7648
rect 13501 7584 13517 7648
rect 13581 7584 13597 7648
rect 13661 7584 13669 7648
rect 13349 6560 13669 7584
rect 13349 6496 13357 6560
rect 13421 6496 13437 6560
rect 13501 6496 13517 6560
rect 13581 6496 13597 6560
rect 13661 6496 13669 6560
rect 13349 5472 13669 6496
rect 13349 5408 13357 5472
rect 13421 5408 13437 5472
rect 13501 5408 13517 5472
rect 13581 5408 13597 5472
rect 13661 5408 13669 5472
rect 13349 4384 13669 5408
rect 13349 4320 13357 4384
rect 13421 4320 13437 4384
rect 13501 4320 13517 4384
rect 13581 4320 13597 4384
rect 13661 4320 13669 4384
rect 13349 3296 13669 4320
rect 13349 3232 13357 3296
rect 13421 3232 13437 3296
rect 13501 3232 13517 3296
rect 13581 3232 13597 3296
rect 13661 3232 13669 3296
rect 13349 2208 13669 3232
rect 13349 2144 13357 2208
rect 13421 2144 13437 2208
rect 13501 2144 13517 2208
rect 13581 2144 13597 2208
rect 13661 2144 13669 2208
rect 13349 1120 13669 2144
rect 13349 1056 13357 1120
rect 13421 1056 13437 1120
rect 13501 1056 13517 1120
rect 13581 1056 13597 1120
rect 13661 1056 13669 1120
rect 13349 496 13669 1056
rect 15200 14720 15520 15280
rect 15200 14656 15208 14720
rect 15272 14656 15288 14720
rect 15352 14656 15368 14720
rect 15432 14656 15448 14720
rect 15512 14656 15520 14720
rect 15200 13632 15520 14656
rect 15200 13568 15208 13632
rect 15272 13568 15288 13632
rect 15352 13568 15368 13632
rect 15432 13568 15448 13632
rect 15512 13568 15520 13632
rect 15200 12544 15520 13568
rect 15200 12480 15208 12544
rect 15272 12480 15288 12544
rect 15352 12480 15368 12544
rect 15432 12480 15448 12544
rect 15512 12480 15520 12544
rect 15200 11456 15520 12480
rect 15200 11392 15208 11456
rect 15272 11392 15288 11456
rect 15352 11392 15368 11456
rect 15432 11392 15448 11456
rect 15512 11392 15520 11456
rect 15200 10368 15520 11392
rect 15200 10304 15208 10368
rect 15272 10304 15288 10368
rect 15352 10304 15368 10368
rect 15432 10304 15448 10368
rect 15512 10304 15520 10368
rect 15200 9280 15520 10304
rect 15200 9216 15208 9280
rect 15272 9216 15288 9280
rect 15352 9216 15368 9280
rect 15432 9216 15448 9280
rect 15512 9216 15520 9280
rect 15200 8192 15520 9216
rect 15200 8128 15208 8192
rect 15272 8128 15288 8192
rect 15352 8128 15368 8192
rect 15432 8128 15448 8192
rect 15512 8128 15520 8192
rect 15200 7104 15520 8128
rect 15200 7040 15208 7104
rect 15272 7040 15288 7104
rect 15352 7040 15368 7104
rect 15432 7040 15448 7104
rect 15512 7040 15520 7104
rect 15200 6016 15520 7040
rect 15200 5952 15208 6016
rect 15272 5952 15288 6016
rect 15352 5952 15368 6016
rect 15432 5952 15448 6016
rect 15512 5952 15520 6016
rect 15200 4928 15520 5952
rect 15200 4864 15208 4928
rect 15272 4864 15288 4928
rect 15352 4864 15368 4928
rect 15432 4864 15448 4928
rect 15512 4864 15520 4928
rect 15200 3840 15520 4864
rect 15200 3776 15208 3840
rect 15272 3776 15288 3840
rect 15352 3776 15368 3840
rect 15432 3776 15448 3840
rect 15512 3776 15520 3840
rect 15200 2752 15520 3776
rect 15200 2688 15208 2752
rect 15272 2688 15288 2752
rect 15352 2688 15368 2752
rect 15432 2688 15448 2752
rect 15512 2688 15520 2752
rect 15200 1664 15520 2688
rect 15200 1600 15208 1664
rect 15272 1600 15288 1664
rect 15352 1600 15368 1664
rect 15432 1600 15448 1664
rect 15512 1600 15520 1664
rect 15200 576 15520 1600
rect 15200 512 15208 576
rect 15272 512 15288 576
rect 15352 512 15368 576
rect 15432 512 15448 576
rect 15512 512 15520 576
rect 15200 496 15520 512
use sky130_fd_sc_hd__xnor2_2  _097_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 10948 0 -1 1632
box -38 -48 1234 592
use sky130_fd_sc_hd__or2b_1  _098_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 12144 0 1 544
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_1  _099_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 11776 0 1 544
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _100_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 12512 0 1 1632
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _101_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 10856 0 1 1632
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _102_
timestamp 1704896540
transform 1 0 11408 0 1 1632
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _103_
timestamp 1704896540
transform 1 0 11132 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _104_
timestamp 1704896540
transform 1 0 10580 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _105_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 11684 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _106_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 11132 0 -1 3808
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _107_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 12052 0 1 2720
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _108_
timestamp 1704896540
transform -1 0 13340 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _109_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 12512 0 -1 2720
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _110_
timestamp 1704896540
transform 1 0 13524 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _111_
timestamp 1704896540
transform 1 0 12420 0 -1 3808
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _112_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 12512 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _113_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 11132 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__and2b_1  _114_
timestamp 1704896540
transform 1 0 10120 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _115_
timestamp 1704896540
transform 1 0 9568 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _116_
timestamp 1704896540
transform 1 0 9936 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _117_
timestamp 1704896540
transform 1 0 11960 0 1 4896
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _118_
timestamp 1704896540
transform 1 0 12604 0 1 4896
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_2  _119_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 14168 0 1 3808
box -38 -48 682 592
use sky130_fd_sc_hd__or3_1  _120_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 12972 0 1 3808
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _121_
timestamp 1704896540
transform -1 0 14628 0 1 3808
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _122_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 13708 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _123_
timestamp 1704896540
transform 1 0 10948 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _124_
timestamp 1704896540
transform 1 0 10304 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _125_
timestamp 1704896540
transform 1 0 11500 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__and3b_1  _126_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 10212 0 -1 4896
box -38 -48 682 592
use sky130_fd_sc_hd__a311o_1  _127_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 11960 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__xor2_1  _128_
timestamp 1704896540
transform 1 0 10948 0 -1 7072
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _129_
timestamp 1704896540
transform -1 0 12236 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _130_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 12236 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  _131_
timestamp 1704896540
transform 1 0 12880 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _132_
timestamp 1704896540
transform 1 0 13524 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _133_
timestamp 1704896540
transform 1 0 13156 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _134_
timestamp 1704896540
transform -1 0 14168 0 1 5984
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _135_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 13524 0 1 7072
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _136_
timestamp 1704896540
transform -1 0 10580 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__xnor2_1  _137_
timestamp 1704896540
transform 1 0 9292 0 1 8160
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _138_
timestamp 1704896540
transform 1 0 11224 0 1 8160
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _139_
timestamp 1704896540
transform 1 0 12052 0 1 8160
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _140_
timestamp 1704896540
transform 1 0 12328 0 -1 8160
box -38 -48 682 592
use sky130_fd_sc_hd__or2b_1  _141_
timestamp 1704896540
transform 1 0 10120 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__or2b_1  _142_
timestamp 1704896540
transform 1 0 9568 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _143_
timestamp 1704896540
transform -1 0 11132 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _144_
timestamp 1704896540
transform 1 0 9384 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _145_
timestamp 1704896540
transform 1 0 10212 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__a2bb2o_1  _146_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 9476 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_1  _147_
timestamp 1704896540
transform -1 0 11224 0 1 8160
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _148_
timestamp 1704896540
transform 1 0 10212 0 1 10336
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _149_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 11592 0 -1 10336
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _150_
timestamp 1704896540
transform 1 0 11316 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _151_
timestamp 1704896540
transform -1 0 12512 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _152_
timestamp 1704896540
transform 1 0 12144 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__a311o_1  _153_
timestamp 1704896540
transform 1 0 12604 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _154_
timestamp 1704896540
transform 1 0 12788 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _155_
timestamp 1704896540
transform 1 0 12788 0 -1 10336
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _156_
timestamp 1704896540
transform 1 0 12328 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__o2bb2a_1  _157_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 12052 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__a21boi_1  _158_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 11500 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _159_
timestamp 1704896540
transform 1 0 9844 0 -1 12512
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _160_
timestamp 1704896540
transform 1 0 10396 0 1 11424
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _161_
timestamp 1704896540
transform 1 0 11408 0 1 11424
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _162_
timestamp 1704896540
transform -1 0 12144 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _163_
timestamp 1704896540
transform 1 0 12880 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _164_
timestamp 1704896540
transform 1 0 12328 0 -1 11424
box -38 -48 682 592
use sky130_fd_sc_hd__o21ba_1  _165_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 12144 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__xnor2_1  _166_
timestamp 1704896540
transform 1 0 11684 0 1 12512
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _167_
timestamp 1704896540
transform 1 0 12696 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _168_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 13248 0 1 544
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _169_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 8648 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _170_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 9660 0 1 1632
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _171_
timestamp 1704896540
transform 1 0 9476 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _172_
timestamp 1704896540
transform 1 0 8372 0 1 1632
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _173_
timestamp 1704896540
transform 1 0 7360 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _174_
timestamp 1704896540
transform 1 0 9200 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _175_
timestamp 1704896540
transform 1 0 9016 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _176_
timestamp 1704896540
transform 1 0 8740 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _177_
timestamp 1704896540
transform 1 0 7268 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _178_
timestamp 1704896540
transform 1 0 9292 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _179_
timestamp 1704896540
transform 1 0 9108 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _180_
timestamp 1704896540
transform 1 0 8556 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _181_
timestamp 1704896540
transform 1 0 7084 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _182_
timestamp 1704896540
transform 1 0 8740 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _183_
timestamp 1704896540
transform 1 0 7360 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _184_
timestamp 1704896540
transform 1 0 9200 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _185_
timestamp 1704896540
transform 1 0 8740 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _186_
timestamp 1704896540
transform 1 0 9568 0 1 544
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _187_
timestamp 1704896540
transform 1 0 9108 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _188_
timestamp 1704896540
transform 1 0 7820 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _189_
timestamp 1704896540
transform 1 0 7176 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _190_
timestamp 1704896540
transform 1 0 7820 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _191_
timestamp 1704896540
transform 1 0 7084 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _192_
timestamp 1704896540
transform 1 0 8372 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _193_
timestamp 1704896540
transform 1 0 7084 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _194_
timestamp 1704896540
transform 1 0 8924 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _195_
timestamp 1704896540
transform 1 0 7452 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _196_
timestamp 1704896540
transform 1 0 8372 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _197_
timestamp 1704896540
transform 1 0 7360 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _198_
timestamp 1704896540
transform 1 0 8372 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _199_
timestamp 1704896540
transform 1 0 7452 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _200_
timestamp 1704896540
transform 1 0 10028 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _201_
timestamp 1704896540
transform -1 0 10396 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__dfstp_1  _202_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 8924 0 -1 2720
box -38 -48 1970 592
use sky130_fd_sc_hd__dfstp_1  _203_
timestamp 1704896540
transform 1 0 6808 0 -1 1632
box -38 -48 1970 592
use sky130_fd_sc_hd__dfstp_1  _204_
timestamp 1704896540
transform 1 0 8556 0 1 3808
box -38 -48 1970 592
use sky130_fd_sc_hd__dfstp_1  _205_
timestamp 1704896540
transform 1 0 6808 0 -1 5984
box -38 -48 1970 592
use sky130_fd_sc_hd__dfstp_1  _206_
timestamp 1704896540
transform 1 0 8740 0 -1 7072
box -38 -48 1970 592
use sky130_fd_sc_hd__dfstp_1  _207_
timestamp 1704896540
transform 1 0 6624 0 -1 9248
box -38 -48 1970 592
use sky130_fd_sc_hd__dfstp_1  _208_
timestamp 1704896540
transform 1 0 6808 0 -1 11424
box -38 -48 1970 592
use sky130_fd_sc_hd__dfstp_1  _209_
timestamp 1704896540
transform 1 0 8188 0 -1 13600
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_4  _210_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 12972 0 -1 1632
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _211_
timestamp 1704896540
transform 1 0 12972 0 -1 2720
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _212_
timestamp 1704896540
transform 1 0 12972 0 -1 3808
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _213_
timestamp 1704896540
transform 1 0 12972 0 -1 5984
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _214_
timestamp 1704896540
transform 1 0 12972 0 -1 8160
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _215_
timestamp 1704896540
transform 1 0 12972 0 -1 9248
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _216_
timestamp 1704896540
transform 1 0 12972 0 -1 11424
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _217_
timestamp 1704896540
transform 1 0 12696 0 -1 12512
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _218_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 8740 0 -1 1632
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _219_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 6348 0 1 2720
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _220_
timestamp 1704896540
transform 1 0 6440 0 1 3808
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _221_
timestamp 1704896540
transform 1 0 6532 0 -1 7072
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _222_
timestamp 1704896540
transform 1 0 6992 0 -1 8160
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _223_
timestamp 1704896540
transform 1 0 6900 0 -1 10336
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _224_
timestamp 1704896540
transform 1 0 6992 0 -1 12512
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _225_
timestamp 1704896540
transform 1 0 10948 0 -1 13600
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_clk $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 11592 0 1 7072
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_0__f_clk
timestamp 1704896540
transform 1 0 9384 0 1 4896
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_1__f_clk
timestamp 1704896540
transform 1 0 9660 0 1 9248
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_4  fanout3
timestamp 1704896540
transform -1 0 8280 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout4
timestamp 1704896540
transform -1 0 9844 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  fanout5 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 9844 0 1 13600
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_3 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 828 0 1 544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_15
timestamp 1704896540
transform 1 0 1932 0 1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_27 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 3036 0 1 544
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_29
timestamp 1704896540
transform 1 0 3220 0 1 544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_41
timestamp 1704896540
transform 1 0 4324 0 1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_53 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 5428 0 1 544
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_57
timestamp 1704896540
transform 1 0 5796 0 1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_69 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 6900 0 1 544
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_73
timestamp 1704896540
transform 1 0 7268 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_0_77 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 7636 0 1 544
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_83
timestamp 1704896540
transform 1 0 8188 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_89
timestamp 1704896540
transform 1 0 8740 0 1 544
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_96 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 9384 0 1 544
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_107
timestamp 1704896540
transform 1 0 10396 0 1 544
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_111
timestamp 1704896540
transform 1 0 10764 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_113 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 10948 0 1 544
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_121
timestamp 1704896540
transform 1 0 11684 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_138
timestamp 1704896540
transform 1 0 13248 0 1 544
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_141
timestamp 1704896540
transform 1 0 13524 0 1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_153
timestamp 1704896540
transform 1 0 14628 0 1 544
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_157
timestamp 1704896540
transform 1 0 14996 0 1 544
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_3
timestamp 1704896540
transform 1 0 828 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_15
timestamp 1704896540
transform 1 0 1932 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_27
timestamp 1704896540
transform 1 0 3036 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_39
timestamp 1704896540
transform 1 0 4140 0 -1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_51
timestamp 1704896540
transform 1 0 5244 0 -1 1632
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_55
timestamp 1704896540
transform 1 0 5612 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1_57
timestamp 1704896540
transform 1 0 5796 0 -1 1632
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1_65
timestamp 1704896540
transform 1 0 6532 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1_109
timestamp 1704896540
transform 1 0 10580 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_134
timestamp 1704896540
transform 1 0 12880 0 -1 1632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_3
timestamp 1704896540
transform 1 0 828 0 1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_15
timestamp 1704896540
transform 1 0 1932 0 1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_27
timestamp 1704896540
transform 1 0 3036 0 1 1632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_29
timestamp 1704896540
transform 1 0 3220 0 1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_41
timestamp 1704896540
transform 1 0 4324 0 1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_53
timestamp 1704896540
transform 1 0 5428 0 1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_65
timestamp 1704896540
transform 1 0 6532 0 1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_77
timestamp 1704896540
transform 1 0 7636 0 1 1632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_83
timestamp 1704896540
transform 1 0 8188 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2_94
timestamp 1704896540
transform 1 0 9200 0 1 1632
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_98
timestamp 1704896540
transform 1 0 9568 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2_108
timestamp 1704896540
transform 1 0 10488 0 1 1632
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_130
timestamp 1704896540
transform 1 0 12512 0 1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_135
timestamp 1704896540
transform 1 0 12972 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_139
timestamp 1704896540
transform 1 0 13340 0 1 1632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_144
timestamp 1704896540
transform 1 0 13800 0 1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_156
timestamp 1704896540
transform 1 0 14904 0 1 1632
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_3
timestamp 1704896540
transform 1 0 828 0 -1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_15
timestamp 1704896540
transform 1 0 1932 0 -1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_27
timestamp 1704896540
transform 1 0 3036 0 -1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_39
timestamp 1704896540
transform 1 0 4140 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_51
timestamp 1704896540
transform 1 0 5244 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_55
timestamp 1704896540
transform 1 0 5612 0 -1 2720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_57
timestamp 1704896540
transform 1 0 5796 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3_69
timestamp 1704896540
transform 1 0 6900 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_75
timestamp 1704896540
transform 1 0 7452 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3_88
timestamp 1704896540
transform 1 0 8648 0 -1 2720
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_113
timestamp 1704896540
transform 1 0 10948 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_125
timestamp 1704896540
transform 1 0 12052 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_129
timestamp 1704896540
transform 1 0 12420 0 -1 2720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_3
timestamp 1704896540
transform 1 0 828 0 1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_15
timestamp 1704896540
transform 1 0 1932 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_27
timestamp 1704896540
transform 1 0 3036 0 1 2720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_29
timestamp 1704896540
transform 1 0 3220 0 1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_41
timestamp 1704896540
transform 1 0 4324 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_4_53
timestamp 1704896540
transform 1 0 5428 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_61
timestamp 1704896540
transform 1 0 6164 0 1 2720
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_85
timestamp 1704896540
transform 1 0 8372 0 1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_100
timestamp 1704896540
transform 1 0 9752 0 1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_112
timestamp 1704896540
transform 1 0 10856 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_124
timestamp 1704896540
transform 1 0 11960 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_4_132
timestamp 1704896540
transform 1 0 12696 0 1 2720
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_141
timestamp 1704896540
transform 1 0 13524 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4_153
timestamp 1704896540
transform 1 0 14628 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_157
timestamp 1704896540
transform 1 0 14996 0 1 2720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_3
timestamp 1704896540
transform 1 0 828 0 -1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_15
timestamp 1704896540
transform 1 0 1932 0 -1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_27
timestamp 1704896540
transform 1 0 3036 0 -1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_39
timestamp 1704896540
transform 1 0 4140 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_51
timestamp 1704896540
transform 1 0 5244 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_55
timestamp 1704896540
transform 1 0 5612 0 -1 3808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_57
timestamp 1704896540
transform 1 0 5796 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_69
timestamp 1704896540
transform 1 0 6900 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_74
timestamp 1704896540
transform 1 0 7360 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_78
timestamp 1704896540
transform 1 0 7728 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_5_103
timestamp 1704896540
transform 1 0 10028 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_111
timestamp 1704896540
transform 1 0 10764 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_113
timestamp 1704896540
transform 1 0 10948 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_122
timestamp 1704896540
transform 1 0 11776 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_128
timestamp 1704896540
transform 1 0 12328 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_134
timestamp 1704896540
transform 1 0 12880 0 -1 3808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_3
timestamp 1704896540
transform 1 0 828 0 1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_15
timestamp 1704896540
transform 1 0 1932 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_27
timestamp 1704896540
transform 1 0 3036 0 1 3808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_29
timestamp 1704896540
transform 1 0 3220 0 1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_41
timestamp 1704896540
transform 1 0 4324 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_6_53
timestamp 1704896540
transform 1 0 5428 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_6_61
timestamp 1704896540
transform 1 0 6164 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_85
timestamp 1704896540
transform 1 0 8372 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_108
timestamp 1704896540
transform 1 0 10488 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_6_124
timestamp 1704896540
transform 1 0 11960 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_6_132
timestamp 1704896540
transform 1 0 12696 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_6_153
timestamp 1704896540
transform 1 0 14628 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_157
timestamp 1704896540
transform 1 0 14996 0 1 3808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_3
timestamp 1704896540
transform 1 0 828 0 -1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_15
timestamp 1704896540
transform 1 0 1932 0 -1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_27
timestamp 1704896540
transform 1 0 3036 0 -1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_39
timestamp 1704896540
transform 1 0 4140 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_51
timestamp 1704896540
transform 1 0 5244 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_55
timestamp 1704896540
transform 1 0 5612 0 -1 4896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_57
timestamp 1704896540
transform 1 0 5796 0 -1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_69
timestamp 1704896540
transform 1 0 6900 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_7_81
timestamp 1704896540
transform 1 0 8004 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_7_89
timestamp 1704896540
transform 1 0 8740 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_95
timestamp 1704896540
transform 1 0 9292 0 -1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_101
timestamp 1704896540
transform 1 0 9844 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_113
timestamp 1704896540
transform 1 0 10948 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_7_119
timestamp 1704896540
transform 1 0 11500 0 -1 4896
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_130
timestamp 1704896540
transform 1 0 12512 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_142
timestamp 1704896540
transform 1 0 13616 0 -1 4896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_146
timestamp 1704896540
transform 1 0 13984 0 -1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_3
timestamp 1704896540
transform 1 0 828 0 1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_15
timestamp 1704896540
transform 1 0 1932 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_27
timestamp 1704896540
transform 1 0 3036 0 1 4896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_29
timestamp 1704896540
transform 1 0 3220 0 1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_41
timestamp 1704896540
transform 1 0 4324 0 1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_53
timestamp 1704896540
transform 1 0 5428 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_8_65
timestamp 1704896540
transform 1 0 6532 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_8_76
timestamp 1704896540
transform 1 0 7544 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_8_85
timestamp 1704896540
transform 1 0 8372 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_8_93
timestamp 1704896540
transform 1 0 9108 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_138
timestamp 1704896540
transform 1 0 13248 0 1 4896
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_144
timestamp 1704896540
transform 1 0 13800 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_156
timestamp 1704896540
transform 1 0 14904 0 1 4896
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_3
timestamp 1704896540
transform 1 0 828 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_15
timestamp 1704896540
transform 1 0 1932 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_27
timestamp 1704896540
transform 1 0 3036 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_39
timestamp 1704896540
transform 1 0 4140 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_51
timestamp 1704896540
transform 1 0 5244 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_55
timestamp 1704896540
transform 1 0 5612 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_9_57
timestamp 1704896540
transform 1 0 5796 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_9_65
timestamp 1704896540
transform 1 0 6532 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_110
timestamp 1704896540
transform 1 0 10672 0 -1 5984
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_113
timestamp 1704896540
transform 1 0 10948 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_9_125
timestamp 1704896540
transform 1 0 12052 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_133
timestamp 1704896540
transform 1 0 12788 0 -1 5984
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_3
timestamp 1704896540
transform 1 0 828 0 1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_15
timestamp 1704896540
transform 1 0 1932 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_27
timestamp 1704896540
transform 1 0 3036 0 1 5984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_29
timestamp 1704896540
transform 1 0 3220 0 1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_41
timestamp 1704896540
transform 1 0 4324 0 1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_53
timestamp 1704896540
transform 1 0 5428 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_65
timestamp 1704896540
transform 1 0 6532 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_10_74
timestamp 1704896540
transform 1 0 7360 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_94
timestamp 1704896540
transform 1 0 9200 0 1 5984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_104
timestamp 1704896540
transform 1 0 10120 0 1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_116
timestamp 1704896540
transform 1 0 11224 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_10_128
timestamp 1704896540
transform 1 0 12328 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_136
timestamp 1704896540
transform 1 0 13064 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_10_148
timestamp 1704896540
transform 1 0 14168 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_156
timestamp 1704896540
transform 1 0 14904 0 1 5984
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_3
timestamp 1704896540
transform 1 0 828 0 -1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_15
timestamp 1704896540
transform 1 0 1932 0 -1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_27
timestamp 1704896540
transform 1 0 3036 0 -1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_39
timestamp 1704896540
transform 1 0 4140 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_51
timestamp 1704896540
transform 1 0 5244 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_55
timestamp 1704896540
transform 1 0 5612 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_11_57
timestamp 1704896540
transform 1 0 5796 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_85
timestamp 1704896540
transform 1 0 8372 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_110
timestamp 1704896540
transform 1 0 10672 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_120
timestamp 1704896540
transform 1 0 11592 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_130
timestamp 1704896540
transform 1 0 12512 0 -1 7072
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_140
timestamp 1704896540
transform 1 0 13432 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_152
timestamp 1704896540
transform 1 0 14536 0 -1 7072
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_3
timestamp 1704896540
transform 1 0 828 0 1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_15
timestamp 1704896540
transform 1 0 1932 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_27
timestamp 1704896540
transform 1 0 3036 0 1 7072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_29
timestamp 1704896540
transform 1 0 3220 0 1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_41
timestamp 1704896540
transform 1 0 4324 0 1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_53
timestamp 1704896540
transform 1 0 5428 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_12_65
timestamp 1704896540
transform 1 0 6532 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_73
timestamp 1704896540
transform 1 0 7268 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_78
timestamp 1704896540
transform 1 0 7728 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_12_85
timestamp 1704896540
transform 1 0 8372 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12_96
timestamp 1704896540
transform 1 0 9384 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_12_120
timestamp 1704896540
transform 1 0 11592 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_12_128
timestamp 1704896540
transform 1 0 12328 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_139
timestamp 1704896540
transform 1 0 13340 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_12_148
timestamp 1704896540
transform 1 0 14168 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_156
timestamp 1704896540
transform 1 0 14904 0 1 7072
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_3
timestamp 1704896540
transform 1 0 828 0 -1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_15
timestamp 1704896540
transform 1 0 1932 0 -1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_27
timestamp 1704896540
transform 1 0 3036 0 -1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_39
timestamp 1704896540
transform 1 0 4140 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_51
timestamp 1704896540
transform 1 0 5244 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_55
timestamp 1704896540
transform 1 0 5612 0 -1 8160
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_57
timestamp 1704896540
transform 1 0 5796 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_69
timestamp 1704896540
transform 1 0 6900 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_100
timestamp 1704896540
transform 1 0 9752 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_122
timestamp 1704896540
transform 1 0 11776 0 -1 8160
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_3
timestamp 1704896540
transform 1 0 828 0 1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_15
timestamp 1704896540
transform 1 0 1932 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_27
timestamp 1704896540
transform 1 0 3036 0 1 8160
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_29
timestamp 1704896540
transform 1 0 3220 0 1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_41
timestamp 1704896540
transform 1 0 4324 0 1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_53
timestamp 1704896540
transform 1 0 5428 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_65
timestamp 1704896540
transform 1 0 6532 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_14_74
timestamp 1704896540
transform 1 0 7360 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_82
timestamp 1704896540
transform 1 0 8096 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_14_85
timestamp 1704896540
transform 1 0 8372 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_93
timestamp 1704896540
transform 1 0 9108 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_14_102
timestamp 1704896540
transform 1 0 9936 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_123
timestamp 1704896540
transform 1 0 11868 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_14_132
timestamp 1704896540
transform 1 0 12696 0 1 8160
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_141
timestamp 1704896540
transform 1 0 13524 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_153
timestamp 1704896540
transform 1 0 14628 0 1 8160
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_3
timestamp 1704896540
transform 1 0 828 0 -1 9248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_15
timestamp 1704896540
transform 1 0 1932 0 -1 9248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_27
timestamp 1704896540
transform 1 0 3036 0 -1 9248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_39
timestamp 1704896540
transform 1 0 4140 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_51
timestamp 1704896540
transform 1 0 5244 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_55
timestamp 1704896540
transform 1 0 5612 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_15_57
timestamp 1704896540
transform 1 0 5796 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_65
timestamp 1704896540
transform 1 0 6532 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_96
timestamp 1704896540
transform 1 0 9384 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_15_109
timestamp 1704896540
transform 1 0 10580 0 -1 9248
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_113
timestamp 1704896540
transform 1 0 10948 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_125
timestamp 1704896540
transform 1 0 12052 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_129
timestamp 1704896540
transform 1 0 12420 0 -1 9248
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_3
timestamp 1704896540
transform 1 0 828 0 1 9248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_15
timestamp 1704896540
transform 1 0 1932 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_27
timestamp 1704896540
transform 1 0 3036 0 1 9248
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_29
timestamp 1704896540
transform 1 0 3220 0 1 9248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_41
timestamp 1704896540
transform 1 0 4324 0 1 9248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_53
timestamp 1704896540
transform 1 0 5428 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_16_65
timestamp 1704896540
transform 1 0 6532 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_73
timestamp 1704896540
transform 1 0 7268 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_16_77
timestamp 1704896540
transform 1 0 7636 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_83
timestamp 1704896540
transform 1 0 8188 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_94
timestamp 1704896540
transform 1 0 9200 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_16_119
timestamp 1704896540
transform 1 0 11500 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_127
timestamp 1704896540
transform 1 0 12236 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_131
timestamp 1704896540
transform 1 0 12604 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_16_136
timestamp 1704896540
transform 1 0 13064 0 1 9248
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_141
timestamp 1704896540
transform 1 0 13524 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_153
timestamp 1704896540
transform 1 0 14628 0 1 9248
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_3
timestamp 1704896540
transform 1 0 828 0 -1 10336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_15
timestamp 1704896540
transform 1 0 1932 0 -1 10336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_27
timestamp 1704896540
transform 1 0 3036 0 -1 10336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_39
timestamp 1704896540
transform 1 0 4140 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_17_51
timestamp 1704896540
transform 1 0 5244 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_55
timestamp 1704896540
transform 1 0 5612 0 -1 10336
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_57
timestamp 1704896540
transform 1 0 5796 0 -1 10336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_89
timestamp 1704896540
transform 1 0 8740 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_17_101
timestamp 1704896540
transform 1 0 9844 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_17_109
timestamp 1704896540
transform 1 0 10580 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_17_113
timestamp 1704896540
transform 1 0 10948 0 -1 10336
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_140
timestamp 1704896540
transform 1 0 13432 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_17_152
timestamp 1704896540
transform 1 0 14536 0 -1 10336
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_3
timestamp 1704896540
transform 1 0 828 0 1 10336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_15
timestamp 1704896540
transform 1 0 1932 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_27
timestamp 1704896540
transform 1 0 3036 0 1 10336
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_29
timestamp 1704896540
transform 1 0 3220 0 1 10336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_41
timestamp 1704896540
transform 1 0 4324 0 1 10336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_53
timestamp 1704896540
transform 1 0 5428 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_18_65
timestamp 1704896540
transform 1 0 6532 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_73
timestamp 1704896540
transform 1 0 7268 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_18_77
timestamp 1704896540
transform 1 0 7636 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_83
timestamp 1704896540
transform 1 0 8188 0 1 10336
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_85
timestamp 1704896540
transform 1 0 8372 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_18_97
timestamp 1704896540
transform 1 0 9476 0 1 10336
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_115
timestamp 1704896540
transform 1 0 11132 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_18_130
timestamp 1704896540
transform 1 0 12512 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_138
timestamp 1704896540
transform 1 0 13248 0 1 10336
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_141
timestamp 1704896540
transform 1 0 13524 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_153
timestamp 1704896540
transform 1 0 14628 0 1 10336
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_3
timestamp 1704896540
transform 1 0 828 0 -1 11424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_15
timestamp 1704896540
transform 1 0 1932 0 -1 11424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_27
timestamp 1704896540
transform 1 0 3036 0 -1 11424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_39
timestamp 1704896540
transform 1 0 4140 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_19_51
timestamp 1704896540
transform 1 0 5244 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_55
timestamp 1704896540
transform 1 0 5612 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_19_57
timestamp 1704896540
transform 1 0 5796 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_19_65
timestamp 1704896540
transform 1 0 6532 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_110
timestamp 1704896540
transform 1 0 10672 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_19_119
timestamp 1704896540
transform 1 0 11500 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_127
timestamp 1704896540
transform 1 0 12236 0 -1 11424
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_3
timestamp 1704896540
transform 1 0 828 0 1 11424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_15
timestamp 1704896540
transform 1 0 1932 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_27
timestamp 1704896540
transform 1 0 3036 0 1 11424
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_29
timestamp 1704896540
transform 1 0 3220 0 1 11424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_41
timestamp 1704896540
transform 1 0 4324 0 1 11424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_53
timestamp 1704896540
transform 1 0 5428 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_20_65
timestamp 1704896540
transform 1 0 6532 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_73
timestamp 1704896540
transform 1 0 7268 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_20_78
timestamp 1704896540
transform 1 0 7728 0 1 11424
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_94
timestamp 1704896540
transform 1 0 9200 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_106
timestamp 1704896540
transform 1 0 10304 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_20_114
timestamp 1704896540
transform 1 0 11040 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_20_137
timestamp 1704896540
transform 1 0 13156 0 1 11424
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_141
timestamp 1704896540
transform 1 0 13524 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_153
timestamp 1704896540
transform 1 0 14628 0 1 11424
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_3
timestamp 1704896540
transform 1 0 828 0 -1 12512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_15
timestamp 1704896540
transform 1 0 1932 0 -1 12512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_27
timestamp 1704896540
transform 1 0 3036 0 -1 12512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_39
timestamp 1704896540
transform 1 0 4140 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_21_51
timestamp 1704896540
transform 1 0 5244 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_55
timestamp 1704896540
transform 1 0 5612 0 -1 12512
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_57
timestamp 1704896540
transform 1 0 5796 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_69
timestamp 1704896540
transform 1 0 6900 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_21_90
timestamp 1704896540
transform 1 0 8832 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_21_98
timestamp 1704896540
transform 1 0 9568 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_21_108
timestamp 1704896540
transform 1 0 10488 0 -1 12512
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_113
timestamp 1704896540
transform 1 0 10948 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_21_125
timestamp 1704896540
transform 1 0 12052 0 -1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_131
timestamp 1704896540
transform 1 0 12604 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_21_155
timestamp 1704896540
transform 1 0 14812 0 -1 12512
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_3
timestamp 1704896540
transform 1 0 828 0 1 12512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_15
timestamp 1704896540
transform 1 0 1932 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_27
timestamp 1704896540
transform 1 0 3036 0 1 12512
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_29
timestamp 1704896540
transform 1 0 3220 0 1 12512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_41
timestamp 1704896540
transform 1 0 4324 0 1 12512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_53
timestamp 1704896540
transform 1 0 5428 0 1 12512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_65
timestamp 1704896540
transform 1 0 6532 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_22_77
timestamp 1704896540
transform 1 0 7636 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_83
timestamp 1704896540
transform 1 0 8188 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_22_85
timestamp 1704896540
transform 1 0 8372 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_92
timestamp 1704896540
transform 1 0 9016 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_22_112
timestamp 1704896540
transform 1 0 10856 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_120
timestamp 1704896540
transform 1 0 11592 0 1 12512
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_128
timestamp 1704896540
transform 1 0 12328 0 1 12512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_141
timestamp 1704896540
transform 1 0 13524 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_153
timestamp 1704896540
transform 1 0 14628 0 1 12512
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_3
timestamp 1704896540
transform 1 0 828 0 -1 13600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_15
timestamp 1704896540
transform 1 0 1932 0 -1 13600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_27
timestamp 1704896540
transform 1 0 3036 0 -1 13600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_39
timestamp 1704896540
transform 1 0 4140 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_23_51
timestamp 1704896540
transform 1 0 5244 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_55
timestamp 1704896540
transform 1 0 5612 0 -1 13600
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_57
timestamp 1704896540
transform 1 0 5796 0 -1 13600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_69
timestamp 1704896540
transform 1 0 6900 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_81
timestamp 1704896540
transform 1 0 8004 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_23_107
timestamp 1704896540
transform 1 0 10396 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_111
timestamp 1704896540
transform 1 0 10764 0 -1 13600
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_141
timestamp 1704896540
transform 1 0 13524 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_153
timestamp 1704896540
transform 1 0 14628 0 -1 13600
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_3
timestamp 1704896540
transform 1 0 828 0 1 13600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_15
timestamp 1704896540
transform 1 0 1932 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_27
timestamp 1704896540
transform 1 0 3036 0 1 13600
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_29
timestamp 1704896540
transform 1 0 3220 0 1 13600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_41
timestamp 1704896540
transform 1 0 4324 0 1 13600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_53
timestamp 1704896540
transform 1 0 5428 0 1 13600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_65
timestamp 1704896540
transform 1 0 6532 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_24_77
timestamp 1704896540
transform 1 0 7636 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_83
timestamp 1704896540
transform 1 0 8188 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_24_85
timestamp 1704896540
transform 1 0 8372 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_93
timestamp 1704896540
transform 1 0 9108 0 1 13600
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_105
timestamp 1704896540
transform 1 0 10212 0 1 13600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_117
timestamp 1704896540
transform 1 0 11316 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_24_129
timestamp 1704896540
transform 1 0 12420 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_24_137
timestamp 1704896540
transform 1 0 13156 0 1 13600
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_141
timestamp 1704896540
transform 1 0 13524 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_24_153
timestamp 1704896540
transform 1 0 14628 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_157
timestamp 1704896540
transform 1 0 14996 0 1 13600
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_3
timestamp 1704896540
transform 1 0 828 0 -1 14688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_15
timestamp 1704896540
transform 1 0 1932 0 -1 14688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_27
timestamp 1704896540
transform 1 0 3036 0 -1 14688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_39
timestamp 1704896540
transform 1 0 4140 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_25_51
timestamp 1704896540
transform 1 0 5244 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_55
timestamp 1704896540
transform 1 0 5612 0 -1 14688
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_57
timestamp 1704896540
transform 1 0 5796 0 -1 14688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_69
timestamp 1704896540
transform 1 0 6900 0 -1 14688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_81
timestamp 1704896540
transform 1 0 8004 0 -1 14688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_93
timestamp 1704896540
transform 1 0 9108 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_25_105
timestamp 1704896540
transform 1 0 10212 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_111
timestamp 1704896540
transform 1 0 10764 0 -1 14688
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_113
timestamp 1704896540
transform 1 0 10948 0 -1 14688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_125
timestamp 1704896540
transform 1 0 12052 0 -1 14688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_137
timestamp 1704896540
transform 1 0 13156 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_25_149
timestamp 1704896540
transform 1 0 14260 0 -1 14688
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_3
timestamp 1704896540
transform 1 0 828 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_26_15
timestamp 1704896540
transform 1 0 1932 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_26
timestamp 1704896540
transform 1 0 2944 0 1 14688
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_29
timestamp 1704896540
transform 1 0 3220 0 1 14688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_41
timestamp 1704896540
transform 1 0 4324 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_26_53
timestamp 1704896540
transform 1 0 5428 0 1 14688
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_57
timestamp 1704896540
transform 1 0 5796 0 1 14688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_69
timestamp 1704896540
transform 1 0 6900 0 1 14688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_85
timestamp 1704896540
transform 1 0 8372 0 1 14688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_97
timestamp 1704896540
transform 1 0 9476 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_26_109
timestamp 1704896540
transform 1 0 10580 0 1 14688
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_113
timestamp 1704896540
transform 1 0 10948 0 1 14688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_125
timestamp 1704896540
transform 1 0 12052 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_26_137
timestamp 1704896540
transform 1 0 13156 0 1 14688
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_141
timestamp 1704896540
transform 1 0 13524 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_26_153
timestamp 1704896540
transform 1 0 14628 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_157
timestamp 1704896540
transform 1 0 14996 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold1 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 13524 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold2
timestamp 1704896540
transform 1 0 12144 0 -1 1632
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  input1
timestamp 1704896540
transform 1 0 8372 0 1 544
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input2
timestamp 1704896540
transform -1 0 8280 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Left_27
timestamp 1704896540
transform 1 0 552 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Right_0
timestamp 1704896540
transform -1 0 15364 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Left_28
timestamp 1704896540
transform 1 0 552 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Right_1
timestamp 1704896540
transform -1 0 15364 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Left_29
timestamp 1704896540
transform 1 0 552 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Right_2
timestamp 1704896540
transform -1 0 15364 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Left_30
timestamp 1704896540
transform 1 0 552 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Right_3
timestamp 1704896540
transform -1 0 15364 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Left_31
timestamp 1704896540
transform 1 0 552 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Right_4
timestamp 1704896540
transform -1 0 15364 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Left_32
timestamp 1704896540
transform 1 0 552 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Right_5
timestamp 1704896540
transform -1 0 15364 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Left_33
timestamp 1704896540
transform 1 0 552 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Right_6
timestamp 1704896540
transform -1 0 15364 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Left_34
timestamp 1704896540
transform 1 0 552 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Right_7
timestamp 1704896540
transform -1 0 15364 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Left_35
timestamp 1704896540
transform 1 0 552 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Right_8
timestamp 1704896540
transform -1 0 15364 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Left_36
timestamp 1704896540
transform 1 0 552 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Right_9
timestamp 1704896540
transform -1 0 15364 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Left_37
timestamp 1704896540
transform 1 0 552 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Right_10
timestamp 1704896540
transform -1 0 15364 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_Left_38
timestamp 1704896540
transform 1 0 552 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_Right_11
timestamp 1704896540
transform -1 0 15364 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_Left_39
timestamp 1704896540
transform 1 0 552 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_Right_12
timestamp 1704896540
transform -1 0 15364 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_13_Left_40
timestamp 1704896540
transform 1 0 552 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_13_Right_13
timestamp 1704896540
transform -1 0 15364 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_14_Left_41
timestamp 1704896540
transform 1 0 552 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_14_Right_14
timestamp 1704896540
transform -1 0 15364 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_15_Left_42
timestamp 1704896540
transform 1 0 552 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_15_Right_15
timestamp 1704896540
transform -1 0 15364 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_16_Left_43
timestamp 1704896540
transform 1 0 552 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_16_Right_16
timestamp 1704896540
transform -1 0 15364 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_17_Left_44
timestamp 1704896540
transform 1 0 552 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_17_Right_17
timestamp 1704896540
transform -1 0 15364 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_18_Left_45
timestamp 1704896540
transform 1 0 552 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_18_Right_18
timestamp 1704896540
transform -1 0 15364 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_19_Left_46
timestamp 1704896540
transform 1 0 552 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_19_Right_19
timestamp 1704896540
transform -1 0 15364 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_20_Left_47
timestamp 1704896540
transform 1 0 552 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_20_Right_20
timestamp 1704896540
transform -1 0 15364 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_21_Left_48
timestamp 1704896540
transform 1 0 552 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_21_Right_21
timestamp 1704896540
transform -1 0 15364 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_22_Left_49
timestamp 1704896540
transform 1 0 552 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_22_Right_22
timestamp 1704896540
transform -1 0 15364 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_23_Left_50
timestamp 1704896540
transform 1 0 552 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_23_Right_23
timestamp 1704896540
transform -1 0 15364 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_24_Left_51
timestamp 1704896540
transform 1 0 552 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_24_Right_24
timestamp 1704896540
transform -1 0 15364 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_25_Left_52
timestamp 1704896540
transform 1 0 552 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_25_Right_25
timestamp 1704896540
transform -1 0 15364 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_26_Left_53
timestamp 1704896540
transform 1 0 552 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_26_Right_26
timestamp 1704896540
transform -1 0 15364 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  sar_control_6 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 14812 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  sar_control_7
timestamp 1704896540
transform 1 0 14812 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  sar_control_8
timestamp 1704896540
transform 1 0 14812 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  sar_control_9
timestamp 1704896540
transform 1 0 14812 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  sar_control_10
timestamp 1704896540
transform 1 0 14812 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  sar_control_11
timestamp 1704896540
transform 1 0 14812 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  sar_control_12
timestamp 1704896540
transform 1 0 14812 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  sar_control_13
timestamp 1704896540
transform 1 0 14812 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  sar_control_14
timestamp 1704896540
transform -1 0 2944 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_54 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 3128 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_55
timestamp 1704896540
transform 1 0 5704 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_56
timestamp 1704896540
transform 1 0 8280 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_57
timestamp 1704896540
transform 1 0 10856 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_58
timestamp 1704896540
transform 1 0 13432 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_59
timestamp 1704896540
transform 1 0 5704 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_60
timestamp 1704896540
transform 1 0 10856 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_61
timestamp 1704896540
transform 1 0 3128 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_62
timestamp 1704896540
transform 1 0 8280 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_63
timestamp 1704896540
transform 1 0 13432 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_64
timestamp 1704896540
transform 1 0 5704 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_65
timestamp 1704896540
transform 1 0 10856 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_66
timestamp 1704896540
transform 1 0 3128 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_67
timestamp 1704896540
transform 1 0 8280 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_68
timestamp 1704896540
transform 1 0 13432 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_69
timestamp 1704896540
transform 1 0 5704 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_70
timestamp 1704896540
transform 1 0 10856 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_71
timestamp 1704896540
transform 1 0 3128 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_72
timestamp 1704896540
transform 1 0 8280 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_73
timestamp 1704896540
transform 1 0 13432 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_74
timestamp 1704896540
transform 1 0 5704 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_75
timestamp 1704896540
transform 1 0 10856 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_76
timestamp 1704896540
transform 1 0 3128 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_77
timestamp 1704896540
transform 1 0 8280 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_78
timestamp 1704896540
transform 1 0 13432 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_79
timestamp 1704896540
transform 1 0 5704 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_80
timestamp 1704896540
transform 1 0 10856 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_81
timestamp 1704896540
transform 1 0 3128 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_82
timestamp 1704896540
transform 1 0 8280 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_83
timestamp 1704896540
transform 1 0 13432 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_84
timestamp 1704896540
transform 1 0 5704 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_85
timestamp 1704896540
transform 1 0 10856 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_86
timestamp 1704896540
transform 1 0 3128 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_87
timestamp 1704896540
transform 1 0 8280 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_88
timestamp 1704896540
transform 1 0 13432 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_89
timestamp 1704896540
transform 1 0 5704 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_90
timestamp 1704896540
transform 1 0 10856 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_91
timestamp 1704896540
transform 1 0 3128 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_92
timestamp 1704896540
transform 1 0 8280 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_93
timestamp 1704896540
transform 1 0 13432 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_94
timestamp 1704896540
transform 1 0 5704 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_95
timestamp 1704896540
transform 1 0 10856 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_96
timestamp 1704896540
transform 1 0 3128 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_97
timestamp 1704896540
transform 1 0 8280 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_98
timestamp 1704896540
transform 1 0 13432 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_99
timestamp 1704896540
transform 1 0 5704 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_100
timestamp 1704896540
transform 1 0 10856 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_101
timestamp 1704896540
transform 1 0 3128 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_102
timestamp 1704896540
transform 1 0 8280 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_103
timestamp 1704896540
transform 1 0 13432 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_104
timestamp 1704896540
transform 1 0 5704 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_105
timestamp 1704896540
transform 1 0 10856 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_106
timestamp 1704896540
transform 1 0 3128 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_107
timestamp 1704896540
transform 1 0 8280 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_108
timestamp 1704896540
transform 1 0 13432 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_109
timestamp 1704896540
transform 1 0 5704 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_110
timestamp 1704896540
transform 1 0 10856 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_111
timestamp 1704896540
transform 1 0 3128 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_112
timestamp 1704896540
transform 1 0 8280 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_113
timestamp 1704896540
transform 1 0 13432 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_114
timestamp 1704896540
transform 1 0 5704 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_115
timestamp 1704896540
transform 1 0 10856 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_116
timestamp 1704896540
transform 1 0 3128 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_117
timestamp 1704896540
transform 1 0 8280 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_118
timestamp 1704896540
transform 1 0 13432 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_119
timestamp 1704896540
transform 1 0 5704 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_120
timestamp 1704896540
transform 1 0 10856 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_121
timestamp 1704896540
transform 1 0 3128 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_122
timestamp 1704896540
transform 1 0 5704 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_123
timestamp 1704896540
transform 1 0 8280 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_124
timestamp 1704896540
transform 1 0 10856 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_125
timestamp 1704896540
transform 1 0 13432 0 1 14688
box -38 -48 130 592
<< labels >>
rlabel metal2 s 8036 14688 8036 14688 4 VGND
rlabel metal1 s 7958 15232 7958 15232 4 VPWR
rlabel metal2 s 9338 2652 9338 2652 4 _000_
rlabel metal1 s 7314 986 7314 986 4 _001_
rlabel metal2 s 8970 4284 8970 4284 4 _002_
rlabel metal1 s 7268 5338 7268 5338 4 _003_
rlabel metal2 s 9154 7004 9154 7004 4 _004_
rlabel metal2 s 7130 8806 7130 8806 4 _005_
rlabel metal1 s 7314 10778 7314 10778 4 _006_
rlabel metal1 s 8694 12954 8694 12954 4 _007_
rlabel metal1 s 9108 986 9108 986 4 _008_
rlabel metal1 s 6946 2618 6946 2618 4 _009_
rlabel metal1 s 6946 3706 6946 3706 4 _010_
rlabel metal1 s 6992 6426 6992 6426 4 _011_
rlabel metal1 s 7406 7514 7406 7514 4 _012_
rlabel metal1 s 7314 9690 7314 9690 4 _013_
rlabel metal1 s 7406 11866 7406 11866 4 _014_
rlabel metal1 s 11270 13464 11270 13464 4 _015_
rlabel metal1 s 11086 11186 11086 11186 4 _016_
rlabel metal2 s 11362 10268 11362 10268 4 _017_
rlabel metal2 s 12006 10336 12006 10336 4 _018_
rlabel metal1 s 12420 9486 12420 9486 4 _019_
rlabel metal1 s 12558 10098 12558 10098 4 _020_
rlabel metal2 s 12558 9316 12558 9316 4 _021_
rlabel metal2 s 12834 8500 12834 8500 4 _022_
rlabel metal2 s 12926 9860 12926 9860 4 _023_
rlabel metal2 s 12282 9962 12282 9962 4 _024_
rlabel metal1 s 12328 11186 12328 11186 4 _025_
rlabel metal2 s 11178 11492 11178 11492 4 _026_
rlabel metal2 s 10534 11934 10534 11934 4 _027_
rlabel metal1 s 11638 11696 11638 11696 4 _028_
rlabel metal1 s 12374 11730 12374 11730 4 _029_
rlabel metal1 s 12650 11628 12650 11628 4 _030_
rlabel metal2 s 12650 11322 12650 11322 4 _031_
rlabel metal1 s 12098 11866 12098 11866 4 _032_
rlabel metal2 s 12834 1360 12834 1360 4 _033_
rlabel metal1 s 9246 3570 9246 3570 4 _034_
rlabel metal1 s 9614 2074 9614 2074 4 _035_
rlabel metal1 s 7636 782 7636 782 4 _036_
rlabel metal2 s 9246 4182 9246 4182 4 _037_
rlabel metal1 s 8188 5134 8188 5134 4 _038_
rlabel metal2 s 9338 6868 9338 6868 4 _039_
rlabel metal1 s 7958 8398 7958 8398 4 _040_
rlabel metal1 s 8188 10574 8188 10574 4 _041_
rlabel metal1 s 9108 12750 9108 12750 4 _042_
rlabel metal1 s 9476 782 9476 782 4 _043_
rlabel metal1 s 7636 2482 7636 2482 4 _044_
rlabel metal1 s 7590 3570 7590 3570 4 _045_
rlabel metal1 s 7866 6222 7866 6222 4 _046_
rlabel metal1 s 8326 7310 8326 7310 4 _047_
rlabel metal1 s 8004 9486 8004 9486 4 _048_
rlabel metal1 s 8050 11662 8050 11662 4 _049_
rlabel metal1 s 10120 12954 10120 12954 4 _050_
rlabel metal1 s 12236 1734 12236 1734 4 _051_
rlabel metal1 s 12006 1836 12006 1836 4 _052_
rlabel metal1 s 12052 986 12052 986 4 _053_
rlabel metal2 s 13110 1326 13110 1326 4 _054_
rlabel metal1 s 11638 1904 11638 1904 4 _055_
rlabel metal2 s 11362 2822 11362 2822 4 _056_
rlabel metal1 s 11914 4080 11914 4080 4 _057_
rlabel metal1 s 11500 4046 11500 4046 4 _058_
rlabel metal1 s 11638 3910 11638 3910 4 _059_
rlabel metal2 s 12374 3298 12374 3298 4 _060_
rlabel metal2 s 12742 2652 12742 2652 4 _061_
rlabel metal1 s 13846 1870 13846 1870 4 _062_
rlabel metal1 s 13570 1904 13570 1904 4 _063_
rlabel metal1 s 13110 4012 13110 4012 4 _064_
rlabel metal2 s 12834 4930 12834 4930 4 _065_
rlabel metal1 s 11684 4522 11684 4522 4 _066_
rlabel metal1 s 10212 4658 10212 4658 4 _067_
rlabel metal1 s 10028 4658 10028 4658 4 _068_
rlabel metal2 s 10718 4896 10718 4896 4 _069_
rlabel metal1 s 12650 5202 12650 5202 4 _070_
rlabel metal1 s 13018 4080 13018 4080 4 _071_
rlabel metal1 s 14490 4012 14490 4012 4 _072_
rlabel metal1 s 14122 4182 14122 4182 4 _073_
rlabel metal1 s 14076 4250 14076 4250 4 _074_
rlabel metal1 s 11730 7888 11730 7888 4 _075_
rlabel metal1 s 10672 8058 10672 8058 4 _076_
rlabel metal2 s 10810 8330 10810 8330 4 _077_
rlabel metal2 s 11362 4964 11362 4964 4 _078_
rlabel metal2 s 10258 8500 10258 8500 4 _079_
rlabel metal1 s 12190 6800 12190 6800 4 _080_
rlabel metal1 s 13294 7344 13294 7344 4 _081_
rlabel metal1 s 12972 7310 12972 7310 4 _082_
rlabel metal2 s 13938 6426 13938 6426 4 _083_
rlabel metal1 s 13570 6222 13570 6222 4 _084_
rlabel metal1 s 13570 6290 13570 6290 4 _085_
rlabel metal1 s 13386 7514 13386 7514 4 _086_
rlabel metal1 s 11454 8466 11454 8466 4 _087_
rlabel metal1 s 10994 8364 10994 8364 4 _088_
rlabel metal2 s 12190 8738 12190 8738 4 _089_
rlabel metal2 s 12650 8058 12650 8058 4 _090_
rlabel metal1 s 10856 11322 10856 11322 4 _091_
rlabel metal1 s 10764 11118 10764 11118 4 _092_
rlabel metal1 s 10442 10540 10442 10540 4 _093_
rlabel metal2 s 9706 9180 9706 9180 4 _094_
rlabel metal1 s 10166 8908 10166 8908 4 _095_
rlabel metal2 s 10718 8636 10718 8636 4 _096_
rlabel metal1 s 12420 7446 12420 7446 4 clk
rlabel metal1 s 9476 5134 9476 5134 4 clknet_0_clk
rlabel metal2 s 13018 3026 13018 3026 4 clknet_1_0__leaf_clk
rlabel metal1 s 12742 12138 12742 12138 4 clknet_1_1__leaf_clk
rlabel metal2 s 7930 0 7986 400 4 comp_in
port 4 nsew
rlabel metal2 s 10534 986 10534 986 4 first\[0\]
rlabel metal1 s 12374 2958 12374 2958 4 first\[1\]
rlabel metal1 s 11086 4114 11086 4114 4 first\[2\]
rlabel metal1 s 10074 5746 10074 5746 4 first\[3\]
rlabel metal2 s 10350 7786 10350 7786 4 first\[4\]
rlabel metal3 s 9798 9027 9798 9027 4 first\[5\]
rlabel metal2 s 8786 11866 8786 11866 4 first\[6\]
rlabel metal1 s 13064 13294 13064 13294 4 first\[7\]
rlabel metal2 s 10166 2108 10166 2108 4 last\[0\]
rlabel metal2 s 11178 1666 11178 1666 4 last\[1\]
rlabel metal1 s 10051 3910 10051 3910 4 last\[2\]
rlabel metal1 s 8947 5814 8947 5814 4 last\[3\]
rlabel metal2 s 10626 7004 10626 7004 4 last\[4\]
rlabel metal2 s 9062 8670 9062 8670 4 last\[5\]
rlabel metal1 s 9614 11118 9614 11118 4 last\[6\]
rlabel metal1 s 9890 12750 9890 12750 4 last\[7\]
rlabel metal1 s 13248 986 13248 986 4 mid\[0\]
rlabel metal1 s 13432 2074 13432 2074 4 mid\[1\]
rlabel metal1 s 13524 4454 13524 4454 4 mid\[2\]
rlabel metal1 s 13432 5814 13432 5814 4 mid\[3\]
rlabel metal1 s 13110 7854 13110 7854 4 mid\[4\]
rlabel metal1 s 13248 9078 13248 9078 4 mid\[5\]
rlabel metal1 s 12926 11288 12926 11288 4 mid\[6\]
rlabel metal1 s 12650 12342 12650 12342 4 mid\[7\]
rlabel metal1 s 8924 3570 8924 3570 4 net1
rlabel metal3 s 15600 11432 16000 11552 4 net10
port 10 nsew
rlabel metal3 s 15372 12308 15372 12308 4 net11
rlabel metal3 s 15372 13124 15372 13124 4 net12
rlabel metal3 s 15372 13940 15372 13940 4 net13
rlabel metal2 s 2714 15419 2714 15419 4 net14
rlabel metal1 s 12374 12750 12374 12750 4 net15
rlabel metal2 s 12742 1020 12742 1020 4 net16
rlabel metal1 s 9062 13838 9062 13838 4 net2
rlabel metal1 s 12006 1462 12006 1462 4 net3
rlabel metal1 s 14122 12233 14122 12233 4 net4
rlabel metal2 s 14030 3094 14030 3094 4 net5
rlabel metal3 s 15600 8168 16000 8288 4 net6
port 6 nsew
rlabel metal3 s 15372 9044 15372 9044 4 net7
rlabel metal3 s 15372 9860 15372 9860 4 net8
rlabel metal3 s 15042 10659 15042 10659 4 net9
rlabel metal2 s 8050 15317 8050 15317 4 reset_in
rlabel metal3 s 10074 1819 10074 1819 4 sar_out[0]
rlabel metal3 s 15042 2499 15042 2499 4 sar_out[1]
rlabel metal2 s 15042 3417 15042 3417 4 sar_out[2]
rlabel metal2 s 9154 5984 9154 5984 4 sar_out[3]
rlabel metal1 s 9338 7854 9338 7854 4 sar_out[4]
rlabel metal2 s 8878 9248 8878 9248 4 sar_out[5]
rlabel metal1 s 14996 11118 14996 11118 4 sar_out[6]
rlabel metal1 s 12650 12682 12650 12682 4 sar_out[7]
flabel metal4 s 15200 496 15520 15280 0 FreeSans 2400 90 0 0 VGND
port 1 nsew
flabel metal4 s 11498 496 11818 15280 0 FreeSans 2400 90 0 0 VGND
port 1 nsew
flabel metal4 s 7796 496 8116 15280 0 FreeSans 2400 90 0 0 VGND
port 1 nsew
flabel metal4 s 4094 496 4414 15280 0 FreeSans 2400 90 0 0 VGND
port 1 nsew
flabel metal4 s 13349 496 13669 15280 0 FreeSans 2400 90 0 0 VPWR
port 2 nsew
flabel metal4 s 9647 496 9967 15280 0 FreeSans 2400 90 0 0 VPWR
port 2 nsew
flabel metal4 s 5945 496 6265 15280 0 FreeSans 2400 90 0 0 VPWR
port 2 nsew
flabel metal4 s 2243 496 2563 15280 0 FreeSans 2400 90 0 0 VPWR
port 2 nsew
flabel metal2 s 13266 15600 13322 16000 0 FreeSans 280 90 0 0 clk
port 3 nsew
flabel metal2 s 7958 200 7958 200 0 FreeSans 280 90 0 0 comp_in
flabel metal2 s 7930 15600 7986 16000 0 FreeSans 280 90 0 0 reset_in
port 5 nsew
flabel metal3 s 15800 8228 15800 8228 0 FreeSans 600 0 0 0 result[0]
flabel metal3 s 15600 8984 16000 9104 0 FreeSans 600 0 0 0 result[1]
port 7 nsew
flabel metal3 s 15600 9800 16000 9920 0 FreeSans 600 0 0 0 result[2]
port 8 nsew
flabel metal3 s 15600 10616 16000 10736 0 FreeSans 600 0 0 0 result[3]
port 9 nsew
flabel metal3 s 15800 11492 15800 11492 0 FreeSans 600 0 0 0 result[4]
flabel metal3 s 15600 12248 16000 12368 0 FreeSans 600 0 0 0 result[5]
port 11 nsew
flabel metal3 s 15600 13064 16000 13184 0 FreeSans 600 0 0 0 result[6]
port 12 nsew
flabel metal3 s 15600 13880 16000 14000 0 FreeSans 600 0 0 0 result[7]
port 13 nsew
flabel metal3 s 15600 1640 16000 1760 0 FreeSans 600 0 0 0 sar_out[0]
port 14 nsew
flabel metal3 s 15600 2456 16000 2576 0 FreeSans 600 0 0 0 sar_out[1]
port 15 nsew
flabel metal3 s 15600 3272 16000 3392 0 FreeSans 600 0 0 0 sar_out[2]
port 16 nsew
flabel metal3 s 15600 4088 16000 4208 0 FreeSans 600 0 0 0 sar_out[3]
port 17 nsew
flabel metal3 s 15600 4904 16000 5024 0 FreeSans 600 0 0 0 sar_out[4]
port 18 nsew
flabel metal3 s 15600 5720 16000 5840 0 FreeSans 600 0 0 0 sar_out[5]
port 19 nsew
flabel metal3 s 15600 6536 16000 6656 0 FreeSans 600 0 0 0 sar_out[6]
port 20 nsew
flabel metal3 s 15600 7352 16000 7472 0 FreeSans 600 0 0 0 sar_out[7]
port 21 nsew
flabel metal2 s 2594 15600 2650 16000 0 FreeSans 280 90 0 0 valid
port 22 nsew
<< properties >>
string FIXED_BBOX 0 0 16000 16000
string GDS_END 660782
string GDS_FILE ../openlane/sar_control/runs/sar_control/results/final/gds/sar_control.gds
string GDS_START 256682
<< end >>
