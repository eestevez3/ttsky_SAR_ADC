magic
tech sky130A
magscale 1 2
timestamp 1757456334
<< error_p >>
rect -29 151 29 157
rect -29 117 -17 151
rect -29 111 29 117
rect -29 -117 29 -111
rect -29 -151 -17 -117
rect -29 -157 29 -151
<< nwell >>
rect -211 -289 211 289
<< pmos >>
rect -15 -70 15 70
<< pdiff >>
rect -73 58 -15 70
rect -73 -58 -61 58
rect -27 -58 -15 58
rect -73 -70 -15 -58
rect 15 58 73 70
rect 15 -58 27 58
rect 61 -58 73 58
rect 15 -70 73 -58
<< pdiffc >>
rect -61 -58 -27 58
rect 27 -58 61 58
<< nsubdiff >>
rect -175 219 -79 253
rect 79 219 175 253
rect -175 157 -141 219
rect 141 157 175 219
rect -175 -219 -141 -157
rect 141 -219 175 -157
rect -175 -253 -79 -219
rect 79 -253 175 -219
<< nsubdiffcont >>
rect -79 219 79 253
rect -175 -157 -141 157
rect 141 -157 175 157
rect -79 -253 79 -219
<< poly >>
rect -33 151 33 167
rect -33 117 -17 151
rect 17 117 33 151
rect -33 101 33 117
rect -15 70 15 101
rect -15 -101 15 -70
rect -33 -117 33 -101
rect -33 -151 -17 -117
rect 17 -151 33 -117
rect -33 -167 33 -151
<< polycont >>
rect -17 117 17 151
rect -17 -151 17 -117
<< locali >>
rect -175 219 -79 253
rect 79 219 175 253
rect -175 157 -141 219
rect 141 157 175 219
rect -33 117 -17 151
rect 17 117 33 151
rect -61 58 -27 74
rect -61 -74 -27 -58
rect 27 58 61 74
rect 27 -74 61 -58
rect -33 -151 -17 -117
rect 17 -151 33 -117
rect -175 -219 -141 -157
rect 141 -219 175 -157
rect -175 -253 -79 -219
rect 79 -253 175 -219
<< viali >>
rect -17 117 17 151
rect -61 -58 -27 58
rect 27 -58 61 58
rect -17 -151 17 -117
<< metal1 >>
rect -29 151 29 157
rect -29 117 -17 151
rect 17 117 29 151
rect -29 111 29 117
rect -67 58 -21 70
rect -67 -58 -61 58
rect -27 -58 -21 58
rect -67 -70 -21 -58
rect 21 58 67 70
rect 21 -58 27 58
rect 61 -58 67 58
rect 21 -70 67 -58
rect -29 -117 29 -111
rect -29 -151 -17 -117
rect 17 -151 29 -117
rect -29 -157 29 -151
<< properties >>
string FIXED_BBOX -158 -236 158 236
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 0.7 l 0.15 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
