magic
tech sky130A
magscale 1 2
timestamp 1755973519
<< pwell >>
rect -201 -1582 201 1582
<< psubdiff >>
rect -165 1512 -69 1546
rect 69 1512 165 1546
rect -165 1450 -131 1512
rect 131 1450 165 1512
rect -165 -1512 -131 -1450
rect 131 -1512 165 -1450
rect -165 -1546 -69 -1512
rect 69 -1546 165 -1512
<< psubdiffcont >>
rect -69 1512 69 1546
rect -165 -1450 -131 1450
rect 131 -1450 165 1450
rect -69 -1546 69 -1512
<< xpolycontact >>
rect -35 984 35 1416
rect -35 -1416 35 -984
<< ppolyres >>
rect -35 -984 35 984
<< locali >>
rect -165 1512 -69 1546
rect 69 1512 165 1546
rect -165 1450 -131 1512
rect 131 1450 165 1512
rect -165 -1512 -131 -1450
rect 131 -1512 165 -1450
rect -165 -1546 -69 -1512
rect 69 -1546 165 -1512
<< viali >>
rect -19 1001 19 1398
rect -19 -1398 19 -1001
<< metal1 >>
rect -25 1398 25 1410
rect -25 1001 -19 1398
rect 19 1001 25 1398
rect -25 989 25 1001
rect -25 -1001 25 -989
rect -25 -1398 -19 -1001
rect 19 -1398 25 -1001
rect -25 -1410 25 -1398
<< properties >>
string FIXED_BBOX -148 -1529 148 1529
string gencell sky130_fd_pr__res_high_po_0p35
string library sky130
string parameters w 0.350 l 10.0 m 1 nx 1 wmin 0.350 lmin 0.50 rho 319.8 val 10.25k dummy 0 dw 0.0 term 194.82 sterm 0.0 caplen 0 guard 1 glc 1 grc 1 gtc 1 gbc 1 compatible {sky130_fd_pr__res_high_po_0p35  sky130_fd_pr__res_high_po_0p69 sky130_fd_pr__res_high_po_1p41  sky130_fd_pr__res_high_po_2p85 sky130_fd_pr__res_high_po_5p73} snake 0 full_metal 1 wmax 0.350 vias 1 n_guard 0 hv_guard 0 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>
