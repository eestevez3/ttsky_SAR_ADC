magic
tech sky130A
magscale 1 2
timestamp 1755275318
<< metal3 >>
rect -386 1652 386 1680
rect -386 1228 302 1652
rect 366 1228 386 1652
rect -386 1200 386 1228
rect -386 932 386 960
rect -386 508 302 932
rect 366 508 386 932
rect -386 480 386 508
rect -386 212 386 240
rect -386 -212 302 212
rect 366 -212 386 212
rect -386 -240 386 -212
rect -386 -508 386 -480
rect -386 -932 302 -508
rect 366 -932 386 -508
rect -386 -960 386 -932
rect -386 -1228 386 -1200
rect -386 -1652 302 -1228
rect 366 -1652 386 -1228
rect -386 -1680 386 -1652
<< via3 >>
rect 302 1228 366 1652
rect 302 508 366 932
rect 302 -212 366 212
rect 302 -932 366 -508
rect 302 -1652 366 -1228
<< mimcap >>
rect -346 1600 54 1640
rect -346 1280 -306 1600
rect 14 1280 54 1600
rect -346 1240 54 1280
rect -346 880 54 920
rect -346 560 -306 880
rect 14 560 54 880
rect -346 520 54 560
rect -346 160 54 200
rect -346 -160 -306 160
rect 14 -160 54 160
rect -346 -200 54 -160
rect -346 -560 54 -520
rect -346 -880 -306 -560
rect 14 -880 54 -560
rect -346 -920 54 -880
rect -346 -1280 54 -1240
rect -346 -1600 -306 -1280
rect 14 -1600 54 -1280
rect -346 -1640 54 -1600
<< mimcapcontact >>
rect -306 1280 14 1600
rect -306 560 14 880
rect -306 -160 14 160
rect -306 -880 14 -560
rect -306 -1600 14 -1280
<< metal4 >>
rect -198 1601 -94 1800
rect 282 1652 386 1800
rect -307 1600 15 1601
rect -307 1280 -306 1600
rect 14 1280 15 1600
rect -307 1279 15 1280
rect -198 881 -94 1279
rect 282 1228 302 1652
rect 366 1228 386 1652
rect 282 932 386 1228
rect -307 880 15 881
rect -307 560 -306 880
rect 14 560 15 880
rect -307 559 15 560
rect -198 161 -94 559
rect 282 508 302 932
rect 366 508 386 932
rect 282 212 386 508
rect -307 160 15 161
rect -307 -160 -306 160
rect 14 -160 15 160
rect -307 -161 15 -160
rect -198 -559 -94 -161
rect 282 -212 302 212
rect 366 -212 386 212
rect 282 -508 386 -212
rect -307 -560 15 -559
rect -307 -880 -306 -560
rect 14 -880 15 -560
rect -307 -881 15 -880
rect -198 -1279 -94 -881
rect 282 -932 302 -508
rect 366 -932 386 -508
rect 282 -1228 386 -932
rect -307 -1280 15 -1279
rect -307 -1600 -306 -1280
rect 14 -1600 15 -1280
rect -307 -1601 15 -1600
rect -198 -1800 -94 -1601
rect 282 -1652 302 -1228
rect 366 -1652 386 -1228
rect 282 -1800 386 -1652
<< properties >>
string FIXED_BBOX -386 1200 94 1680
string gencell sky130_fd_pr__cap_mim_m3_1
string library sky130
string parameters w 2.0 l 2.0 val 9.52 carea 2.00 cperi 0.19 nx 1 ny 5 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1 ccov 100
<< end >>
