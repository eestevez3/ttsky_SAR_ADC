magic
tech sky130A
magscale 1 2
timestamp 1755981703
<< pwell >>
rect 14 3666 86 4264
rect 618 3666 690 4264
rect 1222 3666 1294 4264
rect 1826 3666 1898 4264
rect 2428 3666 2500 4264
rect 3034 3666 3106 4264
<< viali >>
rect -720 -3394 -686 -3234
<< metal1 >>
rect 14 4680 86 4682
rect 618 4680 690 4682
rect 1222 4680 1294 4682
rect -112 4480 88 4680
rect 492 4480 692 4680
rect 1097 4480 1297 4680
rect 1700 4480 1900 4680
rect 2300 4480 2500 4680
rect 2910 4480 3110 4680
rect 3506 4480 3706 4680
rect 4108 4480 4308 4680
rect 14 3666 86 4480
rect 618 3666 690 4480
rect 1222 3666 1294 4480
rect 1826 3666 1898 4480
rect 2428 3666 2500 4480
rect 3034 3666 3106 4480
rect 3632 3666 3704 4480
rect 4235 3666 4307 4480
rect -590 698 -216 768
rect -590 336 -520 698
rect -286 -956 -216 698
rect 14 -956 84 -302
rect 618 -664 688 -302
rect -286 -1026 84 -956
rect 14 -1664 84 -1026
rect 324 -734 688 -664
rect -1000 -3234 -664 -3210
rect -1000 -3394 -720 -3234
rect -686 -3394 -664 -3234
rect -1000 -3410 -664 -3394
rect -1000 -3994 -800 -3864
rect -590 -3994 -520 -3632
rect -1000 -4064 -520 -3994
rect 14 -3994 84 -3632
rect 324 -3994 394 -734
rect 1222 -1232 1292 -302
rect 1826 -664 1896 -302
rect 618 -1302 1292 -1232
rect 618 -1664 688 -1302
rect 1222 -1664 1292 -1302
rect 1525 -734 1896 -664
rect 618 -3994 688 -3632
rect 14 -4064 688 -3994
rect 1222 -3984 1292 -3632
rect 1525 -3984 1595 -734
rect 2430 -1232 2500 -302
rect 3034 -664 3104 -302
rect 1826 -1302 2500 -1232
rect 1826 -1664 1896 -1302
rect 2430 -1664 2500 -1302
rect 2726 -734 3104 -664
rect 1826 -3984 1896 -3632
rect 1222 -4054 1896 -3984
rect 1222 -4064 1292 -4054
rect 1826 -4064 1896 -4054
rect 2430 -3994 2500 -3632
rect 2726 -3994 2796 -734
rect 3632 -1232 3702 -302
rect 3034 -1302 3702 -1232
rect 3034 -1664 3104 -1302
rect 3632 -1664 3702 -1302
rect 4236 -949 4306 -302
rect 4838 -949 5038 -892
rect 4236 -1019 5038 -949
rect 3034 -3994 3104 -3632
rect 2430 -4064 3104 -3994
rect 3632 -3994 3702 -3632
rect 4236 -3994 4306 -1019
rect 4838 -1092 5038 -1019
rect 3632 -4064 4306 -3994
use sky130_fd_pr__res_high_po_0p35_QPS5FG  XR1
timestamp 1755973519
transform 1 0 4271 0 1 1682
box -201 -2582 201 2582
use sky130_fd_pr__res_high_po_0p35_FFK5MY  XR2
timestamp 1755973519
transform 1 0 3667 0 1 -2648
box -201 -1582 201 1582
use sky130_fd_pr__res_high_po_0p35_QPS5FG  XR3
timestamp 1755973519
transform 1 0 3667 0 1 1682
box -201 -2582 201 2582
use sky130_fd_pr__res_high_po_0p35_FFK5MY  XR4
timestamp 1755973519
transform 1 0 3069 0 1 -2648
box -201 -1582 201 1582
use sky130_fd_pr__res_high_po_0p35_QPS5FG  XR5
timestamp 1755973519
transform 1 0 3069 0 1 1682
box -201 -2582 201 2582
use sky130_fd_pr__res_high_po_0p35_FFK5MY  XR6
timestamp 1755973519
transform 1 0 2465 0 1 -2648
box -201 -1582 201 1582
use sky130_fd_pr__res_high_po_0p35_QPS5FG  XR7
timestamp 1755973519
transform 1 0 2465 0 1 1682
box -201 -2582 201 2582
use sky130_fd_pr__res_high_po_0p35_FFK5MY  XR8
timestamp 1755973519
transform 1 0 1861 0 1 -2648
box -201 -1582 201 1582
use sky130_fd_pr__res_high_po_0p35_QPS5FG  XR9
timestamp 1755973519
transform 1 0 1861 0 1 1682
box -201 -2582 201 2582
use sky130_fd_pr__res_high_po_0p35_FFK5MY  XR10
timestamp 1755973519
transform 1 0 1257 0 1 -2648
box -201 -1582 201 1582
use sky130_fd_pr__res_high_po_0p35_QPS5FG  XR11
timestamp 1755973519
transform 1 0 1257 0 1 1682
box -201 -2582 201 2582
use sky130_fd_pr__res_high_po_0p35_FFK5MY  XR12
timestamp 1755973519
transform 1 0 653 0 1 -2648
box -201 -1582 201 1582
use sky130_fd_pr__res_high_po_0p35_QPS5FG  XR13
timestamp 1755973519
transform 1 0 653 0 1 1682
box -201 -2582 201 2582
use sky130_fd_pr__res_high_po_0p35_FFK5MY  XR14
timestamp 1755973519
transform 1 0 49 0 1 -2648
box -201 -1582 201 1582
use sky130_fd_pr__res_high_po_0p35_QPS5FG  XR15
timestamp 1755973519
transform 1 0 49 0 1 1682
box -201 -2582 201 2582
use sky130_fd_pr__res_high_po_0p35_QPS5FG  XR16
timestamp 1755973519
transform 1 0 -555 0 1 -1648
box -201 -2582 201 2582
<< labels >>
flabel metal1 4838 -1092 5038 -892 0 FreeSans 256 0 0 0 dac_out
port 0 nsew
flabel metal1 4108 4480 4308 4680 0 FreeSans 256 0 0 0 b0
port 9 nsew
flabel metal1 1700 4480 1900 4680 0 FreeSans 256 0 0 0 b4
port 4 nsew
flabel metal1 2300 4480 2500 4680 0 FreeSans 256 0 0 0 b3
port 3 nsew
flabel metal1 2910 4480 3110 4680 0 FreeSans 256 0 0 0 b2
port 8 nsew
flabel metal1 3506 4480 3706 4680 0 FreeSans 256 0 0 0 b1
port 2 nsew
flabel metal1 1097 4480 1297 4680 0 FreeSans 256 0 0 0 b5
port 5 nsew
flabel metal1 492 4480 692 4680 0 FreeSans 256 0 0 0 b6
port 7 nsew
flabel metal1 -112 4480 88 4680 0 FreeSans 256 0 0 0 b7
port 6 nsew
flabel metal1 -1000 -4064 -800 -3864 0 FreeSans 256 0 0 0 VSS
port 1 nsew
flabel metal1 -1000 -3410 -800 -3210 0 FreeSans 256 0 0 0 VSUBS
port 10 nsew
<< end >>
