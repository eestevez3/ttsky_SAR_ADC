Simulation of an R2R DAC with Verilator and d_cosim

.lib /home/ttuser/pdk/sky130A/libs.tech/ngspice/sky130.lib.spice tt

* https://sourceforge.net/p/ngspice/ngspice/ci/master/tree/examples/xspice/verilator/

* The digital portion of the circuit is specified in compiled Verilog.
* list the inputs and outputs
adut [ clk reset_in comp_in ] [b7 b6 b5 b4 b3 b2 b1 b0 result7 result6 result5 result4 result3 result2 result1 result0 valid] null dut
.model dut d_cosim simulation="./sar_control.so"


.include "../xschem/simulation/r2r_dac.spice"
.include "../xschem/simulation/Sample_and_Hold.spice"
.include "../xschem/simulation/comparator.spice" 
*.include "../mag/r2r.spice" 

xr2r b0 b1 b2 b3 b4 b5 b6 b7 out 0 0 r2r

* simulate tt output path
R1 out pin_out 500
C1 out 0 5p



**** End of the ADC and its subcircuits.  Begin test circuit ****

.param vcc=1.8
vcc vcc 0 {vcc}

* Digital clock signal

aclock 0 clk clock
.model clock d_osc cntl_array=[-1 1] freq_array=[1Meg 1Meg]

* reset signal

Vreset n_rst 0 PULSE 3 0 1n 20p 20p 1u 500u

.control
tran 100n 400u
plot pin_out
.endc
.end
