** sch_path: /home/ttuser/ttsky_SAR_ADC/xschem/testbench.sch

.include /home/ttuser/pdk/sky130A/libs.ref/sky130_fd_sc_hd/spice/sky130_fd_sc_hd.spice

**.subckt testbench
x1 SH_OUT VSHIN VSS VCC CLK Sample_and_Hold
VCLK CLK VSS pulse(0 1.8 0.2ns 0.2ns 0.2ns 200ns 400ns 200)
VVCC net5 VSS 'VCC'
VVSS VSS 0 0
VIN VSHIN VSS sin(0.4 0.2 3.3MEG)
VVREF VREF VSS 0.9
R1 pin_out1 SH_OUT 5k m=1
C1 SH_OUT VSS .1p m=1
VrSH VCC net5 0
.save i(vrsh)
x2 SH_PARAX_OUT VSHIN VSS VCC CLK Sample_and_Hold_parax
R2 parax_out SH_PARAX_OUT 5k m=1
C2 SH_PARAX_OUT VSS .1p m=1
x3 net1 VSS VB2 VB4 VB5 VB6 VB8 VB7 VB3 VB1 VSS r2r_dac
VB1 VB1 VSS pwl 0n 0 25n 0 25.2n 'VCC' 500n 'VCC' 500.2n 0
R3 dac_out net1 5k m=1
C3 net1 VSS .1p m=1
x4 net2 VSS VB2 VB4 VB5 VB6 VB8 VB7 VB3 VB1 VSS r2r_dac_parax
R4 dac_out2 net2 5k m=1
C4 net2 VSS .01p m=1
R7 test_out net3 5k m=1
C7 net3 VSS .1p m=1
x8 EN_N PLUS MINUS CAL net3 VCC VSS comparator
VB2 PLUS VSS dc 1.8 pwl 0 'VDL'

VCAL r VSS dc 1.8 pwl 0 0 29.9n 0 30.1n 1.8 69.9n 1.8 70.1n 0 219.8n 0 220n 1.8 259.8n 1.8 260n 0
*+749.8n 0 750n 1.8 789.8n 1.8 790n 0 2.25u 0 2.252u 1.8 2.292u 1.8 2.294u 0 3.25u 0 3.252u 1.8 3.292u 1.8 3.294u 0
VEN f VSS dc 1.8 pwl 0 0 29.9n 0 30.1n 1.8 109.9n 1.8 249.8n 1.8 250n 0 750n 0 750.2n 1.8 1.25u 1.8 1.252u 0 1.75u 0 1.752u 1.8
+ 2.25u 1.8 2.252u 0 2.75u 0 2.752u 1.8 3.25u 1.8 3.252u 0 3.75u 0 3.752u 1.8 4.25u 1.8 4.252u 0 4.75u 0 4.752u 1.8
R5 test_out_parax net4 5k m=1
C5 net4 VSS .1p m=1
x5 EN_N PLUS MINUS CAL net4 VCC VSS comparator_parax
VMINUS2 s 0 pwl 0 0.9 70.2n 0.9 70.5n 0.88 109.9n 0.88 110.1n 1.5 170.2n 1.5 170.5n 0.25 209.9n 0.25 210.1n 1.2 250.9n 1.2 251.2n
+ 0.7 280.9n 0.7 281.1n 0.91 310.9n 0.91 311.1n 0.86 451.9n 0.86 452.1n 0.92
VCLK2 clk_in VSS pulse(0 1.8 0.2n 0.2ns 0.2ns 200ns 4us 500)
VRES reset_in VSS pulse(1.8 0 0.2n 0.2ns 0.2ns 200ns 4us 500)
VB4 VB2 VSS pwl 0n 0 50n 0 50.2n 'VCC' 150n 'VCC' 150.2n 0
VB5 VB3 VSS pwl 0n 0 75n 0 75.2n 'VCC' 600n 'VCC' 600.2n 0
VB6 VB4 VSS pwl 0n 0 150n 0 150.2n 'VCC' 600n 'VCC' 600.2n 0
VB3 VB5 VSS pwl 0n 0 250n 0 250.2n 'VCC' 500n 'VCC' 500.2n 0
VB7 VB6 VSS pwl 0n 0 350n 0 350.2n 'VCC' 500n 'VCC' 500.2n 0
VB8 VB7 VSS pwl 0n 0 400n 0 400.2n 'VCC' 500n 'VCC' 500.2n 0
VB9 VB8 VSS pwl 0n 0 450n 0 450.2n 'VCC' 500n 'VCC' 500.2n 0
VMINUS3 MINUS VSS pwl 0 'VDL' 70.2n 'VDL' 250n 'VDL-DELTA' 750n 'VDL-DELTA' 750.2n 'VDL+DELTA' 1.25u 'VDL+DELTA' 1.252u 'VDL-DELTA2'
+ 1.75u 'VDL-DELTA2' 1.752u 'VDL+DELTA2' 2.25u 'VDL+DELTA2' 2.252u 'VDL-DELTA' 2.75u 'VDL-DELTA' 2.752u 'VDL+DELTA' 3.25u 'VDL+DELTA'
+ 3.252u 'VDL-DELTA2' 3.75u 'VDL-DELTA2' 3.752u 'VDL+DELTA2' 4.25u 'VDL+DELTA2' 4.252u 'VDL-DELTA' 4.75u 'VDL-DELTA' 4.752u 'VDL+DELTA2'
+ 5.25u 'VDL+DELTA2'
VCLK1 EN_N VSS pulse(0 1.8 0.2ns 0.2ns 0.2ns 40ns 500ns 200)
VCLK3 CAL VSS pulse(0 1.8 0.2ns 0.2ns 0.2ns 50ns 500ns 200)
**** begin user architecture code

.param mc_mm_switch=1
.param mc_pr_switch=0
.include /home/ttuser/pdk/sky130A/libs.tech/ngspice/corners/tt.spice
.include /home/ttuser/pdk/sky130A/libs.tech/ngspice/r+c/res_typical__cap_typical.spice
.include /home/ttuser/pdk/sky130A/libs.tech/ngspice/r+c/res_typical__cap_typical__lin.spice
.include /home/ttuser/pdk/sky130A/libs.tech/ngspice/corners/tt/specialized_cells.spice



.option chgtol=4e-16 method=gear
.options acct list
.param VCCGAUSS = agauss(1.8, 0.05, 1)
.param VDLGAUSS = agauss(0.9, 0.23, 1)
.param TEMPGAUSS = agauss(40, 30, 1)
.param 'VCC' = 'VCCGAUSS'
.param 'VDL' = 0.1
.param 'DELTA' = 0.002
.param 'DELTA2' = 0.001
.param 'VREF' = 0.9
.option temp = 'TEMPGAUSS'
.option temp = 27
*vvcc VCC 0 1.8
*vvss VSS 0 0
*vvref VREF 0 0.9
*vclk CLK pulse(1ns 1ns 1ns 5ns 10ns 25)
*vvshin VSHIN sin(0.9 0.9 10MEG)


.control
  setseed  8
  reset
  save all
  savecurrents
  op
  write testbench.raw
  reset
  set appendwrite
  *repeat 5
    save all
    tran 1n 5.5u uic
    write testbench.raw
    set appendwrite
    reset
  *end
  quit 0
.endc

**** end user architecture code
**.ends

* expanding   symbol:  Sample_and_Hold.sym # of pins=5
** sym_path: /home/ttuser/ttsky_SAR_ADC/xschem/Sample_and_Hold.sym
** sch_path: /home/ttuser/ttsky_SAR_ADC/xschem/Sample_and_Hold.sch
.subckt Sample_and_Hold SH_OUT SH_IN VSS VCC SH_CLK
*.ipin SH_IN
*.ipin SH_CLK
*.opin SH_OUT
*.ipin VSS
*.ipin VCC
XC1 SH_OUT VSS sky130_fd_pr__cap_mim_m3_1 W=2 L=2 MF=5 m=5
XM6 SH_OUT CLKN SH_IN VCC sky130_fd_pr__pfet_01v8 L=0.15 W=2 nf=2 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM7 SH_IN CLKB SH_OUT VSS sky130_fd_pr__nfet_01v8 L=0.15 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM8 CLKN SH_CLK VSS VSS sky130_fd_pr__nfet_01v8 L=0.15 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM9 CLKN SH_CLK VCC VCC sky130_fd_pr__pfet_01v8 L=0.15 W=2 nf=2 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM10 CLKB CLKN VSS VSS sky130_fd_pr__nfet_01v8 L=0.15 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM1 CLKB CLKN VCC VCC sky130_fd_pr__pfet_01v8 L=0.15 W=2 nf=2 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
.ends


* expanding   symbol:  r2r_dac.sym # of pins=11
** sym_path: /home/ttuser/ttsky_SAR_ADC/xschem/r2r_dac.sym
** sch_path: /home/ttuser/ttsky_SAR_ADC/xschem/r2r_dac.sch
.subckt r2r_dac dac_out VSS b1 b3 b4 b5 b7 b6 b2 b0 VSUBS
*.ipin b0
*.opin dac_out
*.ipin b1
*.ipin b2
*.ipin b3
*.ipin b4
*.ipin b5
*.ipin b6
*.ipin b7
*.ipin VSS
*.ipin VSUBS
XR1 b0 dac_out VSUBS sky130_fd_pr__res_high_po_0p35 L=20 mult=1 m=1
XR2 dac_out net1 VSUBS sky130_fd_pr__res_high_po_0p35 L=10 mult=1 m=1
XR3 b1 net1 VSUBS sky130_fd_pr__res_high_po_0p35 L=20 mult=1 m=1
XR4 net1 net2 VSUBS sky130_fd_pr__res_high_po_0p35 L=10 mult=1 m=1
XR5 b2 net2 VSUBS sky130_fd_pr__res_high_po_0p35 L=20 mult=1 m=1
XR6 net2 net3 VSUBS sky130_fd_pr__res_high_po_0p35 L=10 mult=1 m=1
XR7 b3 net3 VSUBS sky130_fd_pr__res_high_po_0p35 L=20 mult=1 m=1
XR8 net3 net4 VSUBS sky130_fd_pr__res_high_po_0p35 L=10 mult=1 m=1
XR9 b4 net4 VSUBS sky130_fd_pr__res_high_po_0p35 L=20 mult=1 m=1
XR10 net4 net5 VSUBS sky130_fd_pr__res_high_po_0p35 L=10 mult=1 m=1
XR11 b5 net5 VSUBS sky130_fd_pr__res_high_po_0p35 L=20 mult=1 m=1
XR12 net5 net6 VSUBS sky130_fd_pr__res_high_po_0p35 L=10 mult=1 m=1
XR13 b6 net6 VSUBS sky130_fd_pr__res_high_po_0p35 L=20 mult=1 m=1
XR14 net6 net7 VSUBS sky130_fd_pr__res_high_po_0p35 L=10 mult=1 m=1
XR15 b7 net7 VSUBS sky130_fd_pr__res_high_po_0p35 L=20 mult=1 m=1
XR16 net7 VSS VSUBS sky130_fd_pr__res_high_po_0p35 L=20 mult=1 m=1
.ends


* expanding   symbol:  comparator.sym # of pins=7
** sym_path: /home/ttuser/ttsky_SAR_ADC/xschem/comparator.sym
** sch_path: /home/ttuser/ttsky_SAR_ADC/xschem/comparator.sch
.subckt comparator EN_N PLUS MINUS CAL comp_out VCC VSS
*.ipin VCC
*.ipin VSS
*.ipin EN_N
*.ipin PLUS
*.ipin MINUS
*.opin comp_out
*.ipin CAL
v6 net9 VSSI 0
.save i(v6)
XC4 ZERO0 VSS sky130_fd_pr__cap_mim_m3_1 W=4 L=5 MF=1 m=1
XM1 net6 PLUS net7 VSS sky130_fd_pr__nfet_01v8 L=2 W=2 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM2 net5 MINUS net7 VSS sky130_fd_pr__nfet_01v8 L=2 W=2 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM3 net7 VCC VSS VSS sky130_fd_pr__nfet_01v8 L=4 W=2 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM4 net6 net6 VCC VCC sky130_fd_pr__pfet_01v8_lvt L=2 W=2 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM5 net5 net5 VCC VCC sky130_fd_pr__pfet_01v8_lvt L=2 W=2 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM6 net2 PLUS net3 VCC sky130_fd_pr__pfet_01v8 L=2 W=6 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM7 net1 MINUS net3 VCC sky130_fd_pr__pfet_01v8 L=2 W=6 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM8 net2 net2 VSS VSS sky130_fd_pr__nfet_01v8_lvt L=2 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM9 net1 net1 VSS VSS sky130_fd_pr__nfet_01v8_lvt L=2 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM10 net3 VSS VCC VCC sky130_fd_pr__pfet_01v8 L=2 W=1.2 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM14 out2 net8 VCC VCC sky130_fd_pr__pfet_01v8_lvt L=2 W=2 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM11 net8 net6 VSS VSS sky130_fd_pr__nfet_01v8_lvt L=2 W=2 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM12 out2 net5 VSS VSS sky130_fd_pr__nfet_01v8_lvt L=2 W=2 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM13 net8 net8 VCC VCC sky130_fd_pr__pfet_01v8_lvt L=2 W=2 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM15 out1 net4 VSS VSS sky130_fd_pr__nfet_01v8_lvt L=2 W=2 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM16 net4 net4 VSS VSS sky130_fd_pr__nfet_01v8_lvt L=2 W=2 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM17 net4 net1 VCC VCC sky130_fd_pr__pfet_01v8_lvt L=2 W=2 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM18 out1 net2 VCC VCC sky130_fd_pr__pfet_01v8_lvt L=2 W=2 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM19 comp_out out2 VSS VSS sky130_fd_pr__nfet_01v8 L=2 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM20 comp_out out1 VCC VCC sky130_fd_pr__pfet_01v8 L=2 W=2 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM21 comp_out VSS out2 VSS sky130_fd_pr__nfet_01v8 L=7 W=0.7 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM23 comp_out ZERO0 net9 VSS sky130_fd_pr__nfet_01v8_lvt L=3 W=1 nf=1 ad='W * 0.29' as='W * 0.29' pd='2*(W + 0.29)' ps='2*(W + 0.29)'
+ nrd=0 nrs=0 sa=0 sb=0 sd=0 mult=1 m=1
XM24 comp_out ZERO0 VCC VCC sky130_fd_pr__pfet_01v8_lvt L=3 W=3 nf=1 ad='W * 0.29' as='W * 0.29' pd='2*(W + 0.29)' ps='2*(W + 0.29)'
+ nrd=0 nrs=0 sa=0 sb=0 sd=0 mult=1 m=1
XM25 CALB CAL VCC VCC sky130_fd_pr__pfet_01v8 L=0.15 W=2 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM26 CALB CAL VSS VSS sky130_fd_pr__nfet_01v8 L=0.15 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM27 CALBB CALB VSS VSS sky130_fd_pr__nfet_01v8 L=0.15 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM28 CALBB CALB VCC VCC sky130_fd_pr__pfet_01v8 L=0.15 W=2 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM29 VSSI EN_N VSS VSS sky130_fd_pr__nfet_01v8 L=0.15 W=8 nf=1 ad='W * 0.29' as='W * 0.29' pd='W + 2 * 0.29' ps='W + 2 * 0.29' nrd=0
+ nrs=0 sa=0 sb=0 sd=0 mult=2 m=2
XM22 comp_out VSS out1 VSS sky130_fd_pr__nfet_01v8 L=7 W=0.7 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM30 comp_out CALB ZERO0 VCC sky130_fd_pr__pfet_01v8 L=0.15 W=0.7 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM31 comp_out CALBB ZERO0 VSS sky130_fd_pr__nfet_01v8 L=0.15 W=0.42 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
.ends


* expanding   symbol:  Sample_and_Hold_parax.sym # of pins=5
** sym_path: /home/ttuser/ttsky_SAR_ADC/xschem/Sample_and_Hold.sym
.include /home/ttuser/ttsky_SAR_ADC/mag/Sample_and_Hold.sim.spice

* expanding   symbol:  r2r_dac_parax.sym # of pins=11
** sym_path: /home/ttuser/ttsky_SAR_ADC/xschem/r2r_dac.sym
.include /home/ttuser/ttsky_SAR_ADC/mag/r2r_dac.sim.spice

* expanding   symbol:  comparator_parax.sym # of pins=7
** sym_path: /home/ttuser/ttsky_SAR_ADC/xschem/comparator.sym
.include /home/ttuser/ttsky_SAR_ADC/mag/comparator.sim.spice
.end
