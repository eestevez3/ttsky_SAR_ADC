magic
tech sky130A
magscale 1 2
timestamp 1755525365
<< metal1 >>
rect 22550 10104 22950 10110
rect 22950 9704 25202 10104
rect 22550 9698 22950 9704
rect 24517 9125 24699 9131
rect 24699 8943 24869 9125
rect 24517 8937 24869 8943
rect 24687 8629 24869 8937
rect 22969 7147 23029 7153
rect 23029 7087 23507 7147
rect 22969 7081 23029 7087
rect 27002 6370 27182 8180
rect 27002 6184 27182 6190
rect 25608 3260 25788 3266
rect 25788 3080 26312 3260
rect 25608 3074 25788 3080
rect 27874 2072 28054 3524
rect 21356 1562 21362 1962
rect 21762 1562 24278 1962
rect 27868 1892 27874 2072
rect 28054 1892 28060 2072
<< via1 >>
rect 22550 9704 22950 10104
rect 24517 8943 24699 9125
rect 22969 7087 23029 7147
rect 27002 6190 27182 6370
rect 25608 3080 25788 3260
rect 21362 1562 21762 1962
rect 27874 1892 28054 2072
<< metal2 >>
rect 21291 10104 21681 10108
rect 21286 10099 22550 10104
rect 21286 9709 21291 10099
rect 21681 9709 22550 10099
rect 21286 9704 22550 9709
rect 22950 9704 22956 10104
rect 21291 9700 21681 9704
rect 24511 8943 24517 9125
rect 24699 8943 24705 9125
rect 22740 7147 22796 7154
rect 22738 7145 22969 7147
rect 22738 7089 22740 7145
rect 22796 7089 22969 7145
rect 22738 7087 22969 7089
rect 23029 7087 23035 7147
rect 22740 7080 22796 7087
rect 26996 6190 27002 6370
rect 27182 6190 28660 6370
rect 18775 3260 18945 3264
rect 18770 3255 25608 3260
rect 18770 3085 18775 3255
rect 18945 3085 25608 3255
rect 18770 3080 25608 3085
rect 25788 3080 25794 3260
rect 18775 3076 18945 3080
rect 27874 2072 28054 2078
rect 20607 1962 20997 1966
rect 21362 1962 21762 1968
rect 20602 1957 21362 1962
rect 20602 1567 20607 1957
rect 20997 1567 21362 1957
rect 20602 1562 21362 1567
rect 20607 1558 20997 1562
rect 21362 1556 21762 1562
rect 27874 1545 28054 1892
rect 28480 1585 28660 6190
rect 27870 1375 27879 1545
rect 28049 1375 28058 1545
rect 28476 1415 28485 1585
rect 28655 1415 28664 1585
rect 28480 1410 28660 1415
rect 27874 1370 28054 1375
<< via2 >>
rect 21291 9709 21681 10099
rect 24522 8948 24694 9120
rect 22740 7089 22796 7145
rect 18775 3085 18945 3255
rect 20607 1567 20997 1957
rect 27879 1375 28049 1545
rect 28485 1415 28655 1585
<< metal3 >>
rect 28758 44697 28764 44761
rect 28828 44697 28834 44761
rect 28766 14027 28826 44697
rect 22738 13967 28826 14027
rect 16000 10099 21686 10104
rect 16000 9709 21291 10099
rect 21681 9709 21686 10099
rect 16000 9704 21686 9709
rect 201 9024 599 9029
rect 16000 9024 16400 9704
rect 200 9023 16400 9024
rect 200 8625 201 9023
rect 599 8625 16400 9023
rect 200 8624 16400 8625
rect 201 8619 599 8624
rect 22738 7150 22798 13967
rect 24517 9120 24699 9125
rect 24517 8948 24522 9120
rect 24694 8948 24699 9120
rect 22735 7145 22801 7150
rect 22735 7089 22740 7145
rect 22796 7089 22801 7145
rect 22735 7084 22801 7089
rect 24517 3661 24699 8948
rect 18770 3255 18950 3260
rect 18770 3085 18775 3255
rect 18945 3085 18950 3255
rect 18770 633 18950 3085
rect 19853 1962 20251 1967
rect 19852 1961 21002 1962
rect 19852 1563 19853 1961
rect 20251 1957 21002 1961
rect 20251 1567 20607 1957
rect 20997 1567 21002 1957
rect 24518 1717 24698 3661
rect 20251 1563 21002 1567
rect 19852 1562 21002 1563
rect 19853 1557 20251 1562
rect 24513 1539 24519 1717
rect 24697 1539 24703 1717
rect 28480 1585 28660 1590
rect 27874 1545 28054 1550
rect 24518 1538 24698 1539
rect 27874 1375 27879 1545
rect 28049 1375 28054 1545
rect 22635 694 22813 699
rect 27874 694 28054 1375
rect 28480 1415 28485 1585
rect 28655 1415 28660 1585
rect 28480 1205 28660 1415
rect 28475 1027 28481 1205
rect 28659 1027 28665 1205
rect 28480 1026 28660 1027
rect 22634 693 28054 694
rect 18765 455 18771 633
rect 18949 455 18955 633
rect 22634 515 22635 693
rect 22813 515 28054 693
rect 22634 514 28054 515
rect 22635 509 22813 514
rect 18770 454 18950 455
<< via3 >>
rect 28764 44697 28828 44761
rect 201 8625 599 9023
rect 19853 1563 20251 1961
rect 24519 1539 24697 1717
rect 28481 1027 28659 1205
rect 18771 455 18949 633
rect 22635 515 22813 693
<< metal4 >>
rect 6134 44152 6194 45152
rect 6686 44152 6746 45152
rect 7238 44152 7298 45152
rect 7790 44152 7850 45152
rect 8342 44152 8402 45152
rect 8894 44152 8954 45152
rect 9446 44152 9506 45152
rect 9998 44152 10058 45152
rect 10550 44152 10610 45152
rect 11102 44152 11162 45152
rect 11654 44152 11714 45152
rect 12206 44152 12266 45152
rect 12758 44152 12818 45152
rect 13310 44152 13370 45152
rect 13862 44152 13922 45152
rect 14414 44152 14474 45152
rect 14966 44152 15026 45152
rect 15518 44152 15578 45152
rect 16070 44152 16130 45152
rect 16622 44152 16682 45152
rect 17174 44152 17234 45152
rect 17726 44152 17786 45152
rect 18278 44152 18338 45152
rect 18830 44152 18890 45152
rect 19382 44620 19442 45152
rect 19934 44620 19994 45152
rect 20486 44620 20546 45152
rect 21038 44620 21098 45152
rect 21590 44620 21650 45152
rect 22142 44620 22202 45152
rect 22694 44620 22754 45152
rect 23246 44620 23306 45152
rect 23798 44620 23858 45152
rect 24350 44620 24410 45152
rect 24902 44620 24962 45152
rect 25454 44620 25514 45152
rect 26006 44620 26066 45152
rect 26558 44620 26618 45152
rect 27110 44620 27170 45152
rect 27662 44620 27722 45152
rect 28214 44695 28274 45152
rect 28766 44762 28826 45152
rect 28763 44761 28829 44762
rect 28763 44697 28764 44761
rect 28828 44697 28829 44761
rect 28763 44696 28829 44697
rect 29318 44695 29378 45152
rect 200 9023 600 44152
rect 200 8625 201 9023
rect 599 8625 600 9023
rect 200 1000 600 8625
rect 800 43752 19288 44152
rect 800 1962 1200 43752
rect 800 1961 20252 1962
rect 800 1563 19853 1961
rect 20251 1563 20252 1961
rect 800 1562 20252 1563
rect 24518 1717 24698 1718
rect 800 1000 1200 1562
rect 24518 1539 24519 1717
rect 24697 1539 24698 1717
rect 22634 693 22814 694
rect 18770 633 18950 634
rect 18770 455 18771 633
rect 18949 455 18950 633
rect 3314 0 3494 200
rect 7178 0 7358 200
rect 11042 0 11222 200
rect 14906 0 15086 200
rect 18770 0 18950 455
rect 22634 515 22635 693
rect 22813 515 22814 693
rect 22634 0 22814 515
rect 24518 442 24698 1539
rect 28480 1205 28660 1206
rect 28480 1027 28481 1205
rect 28659 1027 28660 1205
rect 24518 262 26678 442
rect 26498 0 26678 262
rect 28480 422 28660 1027
rect 28480 242 30542 422
rect 30362 0 30542 242
use Sample_and_Hold  Sample_and_Hold_0
timestamp 1755345873
transform 1 0 19941 0 1 14010
box 3191 -13206 10548 -1660
<< labels >>
flabel metal4 s 29318 44952 29378 45152 0 FreeSans 480 90 0 0 ena
port 1 nsew signal input
flabel metal4 s 28214 44952 28274 45152 0 FreeSans 480 90 0 0 rst_n
port 2 nsew signal input
flabel metal4 s 30362 0 30542 200 0 FreeSans 960 0 0 0 ua[0]
port 3 nsew signal bidirectional
flabel metal4 s 22634 0 22814 200 0 FreeSans 960 0 0 0 ua[2]
port 5 nsew signal bidirectional
flabel metal4 s 18770 0 18950 200 0 FreeSans 960 0 0 0 ua[3]
port 6 nsew signal bidirectional
flabel metal4 s 14906 0 15086 200 0 FreeSans 960 0 0 0 ua[4]
port 7 nsew signal bidirectional
flabel metal4 s 11042 0 11222 200 0 FreeSans 960 0 0 0 ua[5]
port 8 nsew signal bidirectional
flabel metal4 s 7178 0 7358 200 0 FreeSans 960 0 0 0 ua[6]
port 9 nsew signal bidirectional
flabel metal4 s 3314 0 3494 200 0 FreeSans 960 0 0 0 ua[7]
port 10 nsew signal bidirectional
flabel metal4 s 27662 44952 27722 45152 0 FreeSans 480 90 0 0 ui_in[0]
port 11 nsew signal input
flabel metal4 s 27110 44952 27170 45152 0 FreeSans 480 90 0 0 ui_in[1]
port 12 nsew signal input
flabel metal4 s 26558 44952 26618 45152 0 FreeSans 480 90 0 0 ui_in[2]
port 13 nsew signal input
flabel metal4 s 26006 44952 26066 45152 0 FreeSans 480 90 0 0 ui_in[3]
port 14 nsew signal input
flabel metal4 s 25454 44952 25514 45152 0 FreeSans 480 90 0 0 ui_in[4]
port 15 nsew signal input
flabel metal4 s 24902 44952 24962 45152 0 FreeSans 480 90 0 0 ui_in[5]
port 16 nsew signal input
flabel metal4 s 24350 44952 24410 45152 0 FreeSans 480 90 0 0 ui_in[6]
port 17 nsew signal input
flabel metal4 s 23798 44952 23858 45152 0 FreeSans 480 90 0 0 ui_in[7]
port 18 nsew signal input
flabel metal4 s 23246 44952 23306 45152 0 FreeSans 480 90 0 0 uio_in[0]
port 19 nsew signal input
flabel metal4 s 22694 44952 22754 45152 0 FreeSans 480 90 0 0 uio_in[1]
port 20 nsew signal input
flabel metal4 s 22142 44952 22202 45152 0 FreeSans 480 90 0 0 uio_in[2]
port 21 nsew signal input
flabel metal4 s 21590 44952 21650 45152 0 FreeSans 480 90 0 0 uio_in[3]
port 22 nsew signal input
flabel metal4 s 21038 44952 21098 45152 0 FreeSans 480 90 0 0 uio_in[4]
port 23 nsew signal input
flabel metal4 s 20486 44952 20546 45152 0 FreeSans 480 90 0 0 uio_in[5]
port 24 nsew signal input
flabel metal4 s 19934 44952 19994 45152 0 FreeSans 480 90 0 0 uio_in[6]
port 25 nsew signal input
flabel metal4 s 19382 44952 19442 45152 0 FreeSans 480 90 0 0 uio_in[7]
port 26 nsew signal input
flabel metal4 s 9998 44952 10058 45152 0 FreeSans 480 90 0 0 uio_oe[0]
port 27 nsew signal output
flabel metal4 s 9446 44952 9506 45152 0 FreeSans 480 90 0 0 uio_oe[1]
port 28 nsew signal output
flabel metal4 s 8894 44952 8954 45152 0 FreeSans 480 90 0 0 uio_oe[2]
port 29 nsew signal output
flabel metal4 s 8342 44952 8402 45152 0 FreeSans 480 90 0 0 uio_oe[3]
port 30 nsew signal output
flabel metal4 s 7790 44952 7850 45152 0 FreeSans 480 90 0 0 uio_oe[4]
port 31 nsew signal output
flabel metal4 s 7238 44952 7298 45152 0 FreeSans 480 90 0 0 uio_oe[5]
port 32 nsew signal output
flabel metal4 s 6686 44952 6746 45152 0 FreeSans 480 90 0 0 uio_oe[6]
port 33 nsew signal output
flabel metal4 s 6134 44952 6194 45152 0 FreeSans 480 90 0 0 uio_oe[7]
port 34 nsew signal output
flabel metal4 s 14414 44952 14474 45152 0 FreeSans 480 90 0 0 uio_out[0]
port 35 nsew signal output
flabel metal4 s 13862 44952 13922 45152 0 FreeSans 480 90 0 0 uio_out[1]
port 36 nsew signal output
flabel metal4 s 13310 44952 13370 45152 0 FreeSans 480 90 0 0 uio_out[2]
port 37 nsew signal output
flabel metal4 s 12758 44952 12818 45152 0 FreeSans 480 90 0 0 uio_out[3]
port 38 nsew signal output
flabel metal4 s 12206 44952 12266 45152 0 FreeSans 480 90 0 0 uio_out[4]
port 39 nsew signal output
flabel metal4 s 11654 44952 11714 45152 0 FreeSans 480 90 0 0 uio_out[5]
port 40 nsew signal output
flabel metal4 s 11102 44952 11162 45152 0 FreeSans 480 90 0 0 uio_out[6]
port 41 nsew signal output
flabel metal4 s 10550 44952 10610 45152 0 FreeSans 480 90 0 0 uio_out[7]
port 42 nsew signal output
flabel metal4 s 18830 44952 18890 45152 0 FreeSans 480 90 0 0 uo_out[0]
port 43 nsew signal output
flabel metal4 s 18278 44952 18338 45152 0 FreeSans 480 90 0 0 uo_out[1]
port 44 nsew signal output
flabel metal4 s 17726 44952 17786 45152 0 FreeSans 480 90 0 0 uo_out[2]
port 45 nsew signal output
flabel metal4 s 17174 44952 17234 45152 0 FreeSans 480 90 0 0 uo_out[3]
port 46 nsew signal output
flabel metal4 s 16622 44952 16682 45152 0 FreeSans 480 90 0 0 uo_out[4]
port 47 nsew signal output
flabel metal4 s 16070 44952 16130 45152 0 FreeSans 480 90 0 0 uo_out[5]
port 48 nsew signal output
flabel metal4 s 15518 44952 15578 45152 0 FreeSans 480 90 0 0 uo_out[6]
port 49 nsew signal output
flabel metal4 s 14966 44952 15026 45152 0 FreeSans 480 90 0 0 uo_out[7]
port 50 nsew signal output
flabel metal4 200 1000 600 44152 1 FreeSans 1600 0 0 0 VDPWR
port 51 nsew power bidirectional
flabel metal4 800 1000 1200 44152 1 FreeSans 1600 0 0 0 VGND
port 52 nsew ground bidirectional
flabel metal4 s 26498 0 26678 200 0 FreeSans 960 0 0 0 ua[1]
port 4 nsew signal bidirectional
flabel metal4 s 28766 44952 28826 45152 0 FreeSans 480 90 0 0 clk
port 0 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 32200 45152
<< end >>
