** sch_path: /home/ttuser/ttsky_SAR_ADC/xschem/comparator.sch
.subckt comparator EN_N PLUS MINUS CAL comp_out VCC VSS
*.PININFO VCC:I VSS:I EN_N:I PLUS:I MINUS:I comp_out:O CAL:I
v6 net9 VSSI 0
.save i(v6)
XC4 ZERO0 VSS sky130_fd_pr__cap_mim_m3_1 W=4 L=5 m=1
XM1 net6 PLUS net7 VSS sky130_fd_pr__nfet_01v8 L=2 W=2 nf=1 m=1
XM2 net5 MINUS net7 VSS sky130_fd_pr__nfet_01v8 L=2 W=2 nf=1 m=1
XM3 net7 VCC VSS VSS sky130_fd_pr__nfet_01v8 L=4 W=2 nf=1 m=1
XM4 net6 net6 VCC VCC sky130_fd_pr__pfet_01v8_lvt L=2 W=2 nf=1 m=1
XM5 net5 net5 VCC VCC sky130_fd_pr__pfet_01v8_lvt L=2 W=2 nf=1 m=1
XM6 net2 PLUS net3 VCC sky130_fd_pr__pfet_01v8 L=2 W=6 nf=1 m=1
XM7 net1 MINUS net3 VCC sky130_fd_pr__pfet_01v8 L=2 W=6 nf=1 m=1
XM8 net2 net2 VSS VSS sky130_fd_pr__nfet_01v8_lvt L=2 W=1 nf=1 m=1
XM9 net1 net1 VSS VSS sky130_fd_pr__nfet_01v8_lvt L=2 W=1 nf=1 m=1
XM10 net3 VSS VCC VCC sky130_fd_pr__pfet_01v8 L=2 W=1.2 nf=1 m=1
XM14 out2 net8 VCC VCC sky130_fd_pr__pfet_01v8_lvt L=2 W=2 nf=1 m=1
XM11 net8 net6 VSS VSS sky130_fd_pr__nfet_01v8_lvt L=2 W=2 nf=1 m=1
XM12 out2 net5 VSS VSS sky130_fd_pr__nfet_01v8_lvt L=2 W=2 nf=1 m=1
XM13 net8 net8 VCC VCC sky130_fd_pr__pfet_01v8_lvt L=2 W=2 nf=1 m=1
XM15 out1 net4 VSS VSS sky130_fd_pr__nfet_01v8_lvt L=2 W=2 nf=1 m=1
XM16 net4 net4 VSS VSS sky130_fd_pr__nfet_01v8_lvt L=2 W=2 nf=1 m=1
XM17 net4 net1 VCC VCC sky130_fd_pr__pfet_01v8_lvt L=2 W=2 nf=1 m=1
XM18 out1 net2 VCC VCC sky130_fd_pr__pfet_01v8_lvt L=2 W=2 nf=1 m=1
XM19 comp_out out2 VSS VSS sky130_fd_pr__nfet_01v8 L=2 W=1 nf=1 m=1
XM20 comp_out out1 VCC VCC sky130_fd_pr__pfet_01v8 L=2 W=2 nf=1 m=1
XM21 comp_out VSS out2 VSS sky130_fd_pr__nfet_01v8 L=7 W=0.7 nf=1 m=1
XM23 comp_out ZERO0 net9 VSS sky130_fd_pr__nfet_01v8_lvt L=3 W=1 nf=1 m=1
XM24 comp_out ZERO0 VCC VCC sky130_fd_pr__pfet_01v8_lvt L=3 W=3 nf=1 m=1
XM25 CALB CAL VCC VCC sky130_fd_pr__pfet_01v8 L=0.15 W=2 nf=1 m=1
XM26 CALB CAL VSS VSS sky130_fd_pr__nfet_01v8 L=0.15 W=1 nf=1 m=1
XM27 CALBB CALB VSS VSS sky130_fd_pr__nfet_01v8 L=0.15 W=1 nf=1 m=1
XM28 CALBB CALB VCC VCC sky130_fd_pr__pfet_01v8 L=0.15 W=2 nf=1 m=1
XM29 VSSI EN_N VSS VSS sky130_fd_pr__nfet_01v8 L=0.15 W=8 nf=1 m=2
XM22 comp_out VSS out1 VSS sky130_fd_pr__nfet_01v8 L=7 W=0.7 nf=1 m=1
XM30 comp_out CALB ZERO0 VCC sky130_fd_pr__pfet_01v8 L=0.15 W=0.7 nf=1 m=1
XM31 comp_out CALBB ZERO0 VSS sky130_fd_pr__nfet_01v8 L=0.15 W=0.42 nf=1 m=1
.ends
.end
